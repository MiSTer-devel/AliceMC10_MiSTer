module rom_mc10
(
input clk,
input [12:0] addr,
output [7:0] dout,
input cs );
reg [7:0] q;
always @(posedge clk)
begin
case (addr)
	13'h0: q=8'hF2;
	13'h1: q=8'hBA;
	13'h2: q=8'hF3;
	13'h3: q=8'h35;
	13'h4: q=8'hF2;
	13'h5: q=8'hD5;
	13'h6: q=8'h42;
	13'h7: q=8'h15;
	13'h8: q=8'hF6;
	13'h9: q=8'h2A;
	13'hA: q=8'hF5;
	13'hB: q=8'h4D;
	13'hC: q=8'hF0;
	13'hD: q=8'hB9;
	13'hE: q=8'hF5;
	13'hF: q=8'hC9;
	13'h10: q=8'hF6;
	13'h11: q=8'h8C;
	13'h12: q=8'hF6;
	13'h13: q=8'h86;
	13'h14: q=8'hF6;
	13'h15: q=8'hD2;
	13'h16: q=8'hEF;
	13'h17: q=8'h5F;
	13'h18: q=8'hEE;
	13'h19: q=8'h82;
	13'h1A: q=8'hEC;
	13'h1B: q=8'hED;
	13'h1C: q=8'hEF;
	13'h1D: q=8'h1C;
	13'h1E: q=8'hEE;
	13'h1F: q=8'hA2;
	13'h20: q=8'hEE;
	13'h21: q=8'h8E;
	13'h22: q=8'hEE;
	13'h23: q=8'hAD;
	13'h24: q=8'hEE;
	13'h25: q=8'hC8;
	13'h26: q=8'hEE;
	13'h27: q=8'hCF;
	13'h28: q=8'hFB;
	13'h29: q=8'h9C;
	13'h2A: q=8'hFC;
	13'h2B: q=8'h11;
	13'h2C: q=8'hFB;
	13'h2D: q=8'hED;
	13'h2E: q=8'hEC;
	13'h2F: q=8'hDB;
	13'h30: q=8'h79;
	13'h31: q=8'hEF;
	13'h32: q=8'h80;
	13'h33: q=8'h79;
	13'h34: q=8'hEF;
	13'h35: q=8'h75;
	13'h36: q=8'h7B;
	13'h37: q=8'hF0;
	13'h38: q=8'hF1;
	13'h39: q=8'h7B;
	13'h3A: q=8'hF1;
	13'h3B: q=8'hC8;
	13'h3C: q=8'h7F;
	13'h3D: q=8'hF5;
	13'h3E: q=8'h56;
	13'h3F: q=8'h50;
	13'h40: q=8'hEA;
	13'h41: q=8'h8E;
	13'h42: q=8'h46;
	13'h43: q=8'hEA;
	13'h44: q=8'h8D;
	13'h45: q=8'h46;
	13'h46: q=8'h4F;
	13'h47: q=8'hD2;
	13'h48: q=8'h47;
	13'h49: q=8'h4F;
	13'h4A: q=8'h54;
	13'h4B: q=8'hCF;
	13'h4C: q=8'h47;
	13'h4D: q=8'h4F;
	13'h4E: q=8'h53;
	13'h4F: q=8'h55;
	13'h50: q=8'hC2;
	13'h51: q=8'h52;
	13'h52: q=8'h45;
	13'h53: q=8'hCD;
	13'h54: q=8'h49;
	13'h55: q=8'hC6;
	13'h56: q=8'h44;
	13'h57: q=8'h41;
	13'h58: q=8'h54;
	13'h59: q=8'hC1;
	13'h5A: q=8'h50;
	13'h5B: q=8'h52;
	13'h5C: q=8'h49;
	13'h5D: q=8'h4E;
	13'h5E: q=8'hD4;
	13'h5F: q=8'h4F;
	13'h60: q=8'hCE;
	13'h61: q=8'h49;
	13'h62: q=8'h4E;
	13'h63: q=8'h50;
	13'h64: q=8'h55;
	13'h65: q=8'hD4;
	13'h66: q=8'h45;
	13'h67: q=8'h4E;
	13'h68: q=8'hC4;
	13'h69: q=8'h4E;
	13'h6A: q=8'h45;
	13'h6B: q=8'h58;
	13'h6C: q=8'hD4;
	13'h6D: q=8'h44;
	13'h6E: q=8'h49;
	13'h6F: q=8'hCD;
	13'h70: q=8'h52;
	13'h71: q=8'h45;
	13'h72: q=8'h41;
	13'h73: q=8'hC4;
	13'h74: q=8'h4C;
	13'h75: q=8'h45;
	13'h76: q=8'hD4;
	13'h77: q=8'h52;
	13'h78: q=8'h55;
	13'h79: q=8'hCE;
	13'h7A: q=8'h52;
	13'h7B: q=8'h45;
	13'h7C: q=8'h53;
	13'h7D: q=8'h54;
	13'h7E: q=8'h4F;
	13'h7F: q=8'h52;
	13'h80: q=8'hC5;
	13'h81: q=8'h52;
	13'h82: q=8'h45;
	13'h83: q=8'h54;
	13'h84: q=8'h55;
	13'h85: q=8'h52;
	13'h86: q=8'hCE;
	13'h87: q=8'h53;
	13'h88: q=8'h54;
	13'h89: q=8'h4F;
	13'h8A: q=8'hD0;
	13'h8B: q=8'h50;
	13'h8C: q=8'h4F;
	13'h8D: q=8'h4B;
	13'h8E: q=8'hC5;
	13'h8F: q=8'h43;
	13'h90: q=8'h4F;
	13'h91: q=8'h4E;
	13'h92: q=8'hD4;
	13'h93: q=8'h4C;
	13'h94: q=8'h49;
	13'h95: q=8'h53;
	13'h96: q=8'hD4;
	13'h97: q=8'h43;
	13'h98: q=8'h4C;
	13'h99: q=8'h45;
	13'h9A: q=8'h41;
	13'h9B: q=8'hD2;
	13'h9C: q=8'h4E;
	13'h9D: q=8'h45;
	13'h9E: q=8'hD7;
	13'h9F: q=8'h43;
	13'hA0: q=8'h4C;
	13'hA1: q=8'h4F;
	13'hA2: q=8'h41;
	13'hA3: q=8'hC4;
	13'hA4: q=8'h43;
	13'hA5: q=8'h53;
	13'hA6: q=8'h41;
	13'hA7: q=8'h56;
	13'hA8: q=8'hC5;
	13'hA9: q=8'h4C;
	13'hAA: q=8'h4C;
	13'hAB: q=8'h49;
	13'hAC: q=8'h53;
	13'hAD: q=8'hD4;
	13'hAE: q=8'h4C;
	13'hAF: q=8'h50;
	13'hB0: q=8'h52;
	13'hB1: q=8'h49;
	13'hB2: q=8'h4E;
	13'hB3: q=8'hD4;
	13'hB4: q=8'h53;
	13'hB5: q=8'h45;
	13'hB6: q=8'hD4;
	13'hB7: q=8'h52;
	13'hB8: q=8'h45;
	13'hB9: q=8'h53;
	13'hBA: q=8'h45;
	13'hBB: q=8'hD4;
	13'hBC: q=8'h43;
	13'hBD: q=8'h4C;
	13'hBE: q=8'hD3;
	13'hBF: q=8'h53;
	13'hC0: q=8'h4F;
	13'hC1: q=8'h55;
	13'hC2: q=8'h4E;
	13'hC3: q=8'hC4;
	13'hC4: q=8'h45;
	13'hC5: q=8'h58;
	13'hC6: q=8'h45;
	13'hC7: q=8'hC3;
	13'hC8: q=8'h53;
	13'hC9: q=8'h4B;
	13'hCA: q=8'h49;
	13'hCB: q=8'h50;
	13'hCC: q=8'hC6;
	13'hCD: q=8'h54;
	13'hCE: q=8'h41;
	13'hCF: q=8'h42;
	13'hD0: q=8'hA8;
	13'hD1: q=8'h54;
	13'hD2: q=8'hCF;
	13'hD3: q=8'h54;
	13'hD4: q=8'h48;
	13'hD5: q=8'h45;
	13'hD6: q=8'hCE;
	13'hD7: q=8'h4E;
	13'hD8: q=8'h4F;
	13'hD9: q=8'hD4;
	13'hDA: q=8'h53;
	13'hDB: q=8'h54;
	13'hDC: q=8'h45;
	13'hDD: q=8'hD0;
	13'hDE: q=8'h4F;
	13'hDF: q=8'h46;
	13'hE0: q=8'hC6;
	13'hE1: q=8'hAB;
	13'hE2: q=8'hAD;
	13'hE3: q=8'hAA;
	13'hE4: q=8'hAF;
	13'hE5: q=8'hDE;
	13'hE6: q=8'h41;
	13'hE7: q=8'h4E;
	13'hE8: q=8'hC4;
	13'hE9: q=8'h4F;
	13'hEA: q=8'hD2;
	13'hEB: q=8'hBE;
	13'hEC: q=8'hBD;
	13'hED: q=8'hBC;
	13'hEE: q=8'h53;
	13'hEF: q=8'h47;
	13'hF0: q=8'hCE;
	13'hF1: q=8'h49;
	13'hF2: q=8'h4E;
	13'hF3: q=8'hD4;
	13'hF4: q=8'h41;
	13'hF5: q=8'h42;
	13'hF6: q=8'hD3;
	13'hF7: q=8'h55;
	13'hF8: q=8'h53;
	13'hF9: q=8'hD2;
	13'hFA: q=8'h52;
	13'hFB: q=8'h4E;
	13'hFC: q=8'hC4;
	13'hFD: q=8'h53;
	13'hFE: q=8'h51;
	13'hFF: q=8'hD2;
	13'h100: q=8'h4C;
	13'h101: q=8'h4F;
	13'h102: q=8'hC7;
	13'h103: q=8'h45;
	13'h104: q=8'h58;
	13'h105: q=8'hD0;
	13'h106: q=8'h53;
	13'h107: q=8'h49;
	13'h108: q=8'hCE;
	13'h109: q=8'h43;
	13'h10A: q=8'h4F;
	13'h10B: q=8'hD3;
	13'h10C: q=8'h54;
	13'h10D: q=8'h41;
	13'h10E: q=8'hCE;
	13'h10F: q=8'h50;
	13'h110: q=8'h45;
	13'h111: q=8'h45;
	13'h112: q=8'hCB;
	13'h113: q=8'h4C;
	13'h114: q=8'h45;
	13'h115: q=8'hCE;
	13'h116: q=8'h53;
	13'h117: q=8'h54;
	13'h118: q=8'h52;
	13'h119: q=8'hA4;
	13'h11A: q=8'h56;
	13'h11B: q=8'h41;
	13'h11C: q=8'hCC;
	13'h11D: q=8'h41;
	13'h11E: q=8'h53;
	13'h11F: q=8'hC3;
	13'h120: q=8'h43;
	13'h121: q=8'h48;
	13'h122: q=8'h52;
	13'h123: q=8'hA4;
	13'h124: q=8'h4C;
	13'h125: q=8'h45;
	13'h126: q=8'h46;
	13'h127: q=8'h54;
	13'h128: q=8'hA4;
	13'h129: q=8'h52;
	13'h12A: q=8'h49;
	13'h12B: q=8'h47;
	13'h12C: q=8'h48;
	13'h12D: q=8'h54;
	13'h12E: q=8'hA4;
	13'h12F: q=8'h4D;
	13'h130: q=8'h49;
	13'h131: q=8'h44;
	13'h132: q=8'hA4;
	13'h133: q=8'h50;
	13'h134: q=8'h4F;
	13'h135: q=8'h49;
	13'h136: q=8'h4E;
	13'h137: q=8'hD4;
	13'h138: q=8'h56;
	13'h139: q=8'h41;
	13'h13A: q=8'h52;
	13'h13B: q=8'h50;
	13'h13C: q=8'h54;
	13'h13D: q=8'hD2;
	13'h13E: q=8'h49;
	13'h13F: q=8'h4E;
	13'h140: q=8'h4B;
	13'h141: q=8'h45;
	13'h142: q=8'h59;
	13'h143: q=8'hA4;
	13'h144: q=8'h4D;
	13'h145: q=8'h45;
	13'h146: q=8'hCD;
	13'h147: q=8'h0;
	13'h148: q=8'hE4;
	13'h149: q=8'hC4;
	13'h14A: q=8'hE6;
	13'h14B: q=8'h1A;
	13'h14C: q=8'hE6;
	13'h14D: q=8'h4;
	13'h14E: q=8'hE6;
	13'h14F: q=8'h85;
	13'h150: q=8'hE6;
	13'h151: q=8'h72;
	13'h152: q=8'hE6;
	13'h153: q=8'h51;
	13'h154: q=8'hE7;
	13'h155: q=8'h1F;
	13'h156: q=8'hE6;
	13'h157: q=8'h92;
	13'h158: q=8'hE7;
	13'h159: q=8'hDE;
	13'h15A: q=8'hE5;
	13'h15B: q=8'h7F;
	13'h15C: q=8'hE8;
	13'h15D: q=8'hBB;
	13'h15E: q=8'hEB;
	13'h15F: q=8'h12;
	13'h160: q=8'hE8;
	13'h161: q=8'hE;
	13'h162: q=8'hE6;
	13'h163: q=8'hD3;
	13'h164: q=8'hE5;
	13'h165: q=8'hFA;
	13'h166: q=8'hE5;
	13'h167: q=8'h60;
	13'h168: q=8'hE6;
	13'h169: q=8'h31;
	13'h16A: q=8'hE5;
	13'h16B: q=8'h7E;
	13'h16C: q=8'hEF;
	13'h16D: q=8'h66;
	13'h16E: q=8'hE5;
	13'h16F: q=8'hA6;
	13'h170: q=8'hE4;
	13'h171: q=8'hD;
	13'h172: q=8'hE5;
	13'h173: q=8'hB8;
	13'h174: q=8'hE3;
	13'h175: q=8'hCD;
	13'h176: q=8'hFD;
	13'h177: q=8'h5C;
	13'h178: q=8'hFC;
	13'h179: q=8'h3B;
	13'h17A: q=8'hE4;
	13'h17B: q=8'hB;
	13'h17C: q=8'hE7;
	13'h17D: q=8'h1C;
	13'h17E: q=8'hFB;
	13'h17F: q=8'h25;
	13'h180: q=8'hFB;
	13'h181: q=8'h55;
	13'h182: q=8'hFB;
	13'h183: q=8'hBF;
	13'h184: q=8'hFF;
	13'h185: q=8'hA5;
	13'h186: q=8'hFC;
	13'h187: q=8'h4;
	13'h188: q=8'hFE;
	13'h189: q=8'h2F;
	13'h18A: q=8'h4E;
	13'h18B: q=8'h46;
	13'h18C: q=8'h53;
	13'h18D: q=8'h4E;
	13'h18E: q=8'h52;
	13'h18F: q=8'h47;
	13'h190: q=8'h4F;
	13'h191: q=8'h44;
	13'h192: q=8'h46;
	13'h193: q=8'h43;
	13'h194: q=8'h4F;
	13'h195: q=8'h56;
	13'h196: q=8'h4F;
	13'h197: q=8'h4D;
	13'h198: q=8'h55;
	13'h199: q=8'h4C;
	13'h19A: q=8'h42;
	13'h19B: q=8'h53;
	13'h19C: q=8'h44;
	13'h19D: q=8'h44;
	13'h19E: q=8'h2F;
	13'h19F: q=8'h30;
	13'h1A0: q=8'h49;
	13'h1A1: q=8'h44;
	13'h1A2: q=8'h54;
	13'h1A3: q=8'h4D;
	13'h1A4: q=8'h4F;
	13'h1A5: q=8'h53;
	13'h1A6: q=8'h4C;
	13'h1A7: q=8'h53;
	13'h1A8: q=8'h53;
	13'h1A9: q=8'h54;
	13'h1AA: q=8'h43;
	13'h1AB: q=8'h4E;
	13'h1AC: q=8'h49;
	13'h1AD: q=8'h4F;
	13'h1AE: q=8'h46;
	13'h1AF: q=8'h4D;
	13'h1B0: q=8'h20;
	13'h1B1: q=8'h45;
	13'h1B2: q=8'h52;
	13'h1B3: q=8'h52;
	13'h1B4: q=8'h4F;
	13'h1B5: q=8'h52;
	13'h1B6: q=8'h0;
	13'h1B7: q=8'h20;
	13'h1B8: q=8'h49;
	13'h1B9: q=8'h4E;
	13'h1BA: q=8'h20;
	13'h1BB: q=8'h0;
	13'h1BC: q=8'hD;
	13'h1BD: q=8'h4F;
	13'h1BE: q=8'h4B;
	13'h1BF: q=8'hD;
	13'h1C0: q=8'h0;
	13'h1C1: q=8'hD;
	13'h1C2: q=8'h42;
	13'h1C3: q=8'h52;
	13'h1C4: q=8'h45;
	13'h1C5: q=8'h41;
	13'h1C6: q=8'h4B;
	13'h1C7: q=8'h0;
	13'h1C8: q=8'h81;
	13'h1C9: q=8'h3A;
	13'h1CA: q=8'h24;
	13'h1CB: q=8'hB;
	13'h1CC: q=8'h81;
	13'h1CD: q=8'h20;
	13'h1CE: q=8'h26;
	13'h1CF: q=8'h3;
	13'h1D0: q=8'h7E;
	13'h1D1: q=8'h0;
	13'h1D2: q=8'hEB;
	13'h1D3: q=8'h80;
	13'h1D4: q=8'h30;
	13'h1D5: q=8'h80;
	13'h1D6: q=8'hD0;
	13'h1D7: q=8'h39;
	13'h1D8: q=8'h30;
	13'h1D9: q=8'hC6;
	13'h1DA: q=8'h4;
	13'h1DB: q=8'h3A;
	13'h1DC: q=8'hC6;
	13'h1DD: q=8'h12;
	13'h1DE: q=8'hDF;
	13'h1DF: q=8'h89;
	13'h1E0: q=8'hA6;
	13'h1E1: q=8'h0;
	13'h1E2: q=8'h80;
	13'h1E3: q=8'h80;
	13'h1E4: q=8'h26;
	13'h1E5: q=8'h14;
	13'h1E6: q=8'hEE;
	13'h1E7: q=8'h1;
	13'h1E8: q=8'hDF;
	13'h1E9: q=8'h8B;
	13'h1EA: q=8'hDE;
	13'h1EB: q=8'hB5;
	13'h1EC: q=8'h27;
	13'h1ED: q=8'h8;
	13'h1EE: q=8'h9C;
	13'h1EF: q=8'h8B;
	13'h1F0: q=8'h27;
	13'h1F1: q=8'h8;
	13'h1F2: q=8'h8D;
	13'h1F3: q=8'h3B;
	13'h1F4: q=8'h20;
	13'h1F5: q=8'hE6;
	13'h1F6: q=8'hDE;
	13'h1F7: q=8'h8B;
	13'h1F8: q=8'hDF;
	13'h1F9: q=8'hB5;
	13'h1FA: q=8'hDE;
	13'h1FB: q=8'h89;
	13'h1FC: q=8'h4D;
	13'h1FD: q=8'h39;
	13'h1FE: q=8'h8D;
	13'h1FF: q=8'h1E;
	13'h200: q=8'h7;
	13'h201: q=8'h36;
	13'h202: q=8'h9F;
	13'h203: q=8'h91;
	13'h204: q=8'hF;
	13'h205: q=8'h9E;
	13'h206: q=8'hBB;
	13'h207: q=8'hDE;
	13'h208: q=8'hBD;
	13'h209: q=8'h8;
	13'h20A: q=8'h9;
	13'h20B: q=8'hA6;
	13'h20C: q=8'h0;
	13'h20D: q=8'h36;
	13'h20E: q=8'h9C;
	13'h20F: q=8'hC1;
	13'h210: q=8'h26;
	13'h211: q=8'hF8;
	13'h212: q=8'h31;
	13'h213: q=8'h9F;
	13'h214: q=8'hBF;
	13'h215: q=8'h9E;
	13'h216: q=8'h91;
	13'h217: q=8'h32;
	13'h218: q=8'h6;
	13'h219: q=8'h39;
	13'h21A: q=8'h4F;
	13'h21B: q=8'h58;
	13'h21C: q=8'hD3;
	13'h21D: q=8'h99;
	13'h21E: q=8'hC3;
	13'h21F: q=8'h0;
	13'h220: q=8'h3A;
	13'h221: q=8'h25;
	13'h222: q=8'h13;
	13'h223: q=8'h9F;
	13'h224: q=8'h91;
	13'h225: q=8'h93;
	13'h226: q=8'h91;
	13'h227: q=8'h24;
	13'h228: q=8'hD;
	13'h229: q=8'hD3;
	13'h22A: q=8'h91;
	13'h22B: q=8'h39;
	13'h22C: q=8'h4F;
	13'h22D: q=8'hDF;
	13'h22E: q=8'h89;
	13'h22F: q=8'hD3;
	13'h230: q=8'h89;
	13'h231: q=8'hDD;
	13'h232: q=8'h8B;
	13'h233: q=8'hDE;
	13'h234: q=8'h8B;
	13'h235: q=8'h39;
	13'h236: q=8'hC6;
	13'h237: q=8'hC;
	13'h238: q=8'hBD;
	13'h239: q=8'h42;
	13'h23A: q=8'h97;
	13'h23B: q=8'hBD;
	13'h23C: q=8'h42;
	13'h23D: q=8'h9A;
	13'h23E: q=8'hBD;
	13'h23F: q=8'hFC;
	13'h240: q=8'h86;
	13'h241: q=8'hB6;
	13'h242: q=8'h42;
	13'h243: q=8'h6E;
	13'h244: q=8'h27;
	13'h245: q=8'h3;
	13'h246: q=8'hBD;
	13'h247: q=8'hE3;
	13'h248: q=8'hCF;
	13'h249: q=8'hBD;
	13'h24A: q=8'hE3;
	13'h24B: q=8'hEE;
	13'h24C: q=8'h7F;
	13'h24D: q=8'h0;
	13'h24E: q=8'hE8;
	13'h24F: q=8'hBD;
	13'h250: q=8'hE7;
	13'h251: q=8'h6A;
	13'h252: q=8'hBD;
	13'h253: q=8'hE7;
	13'h254: q=8'hBC;
	13'h255: q=8'hCE;
	13'h256: q=8'hE1;
	13'h257: q=8'h8A;
	13'h258: q=8'h3A;
	13'h259: q=8'hA6;
	13'h25A: q=8'h0;
	13'h25B: q=8'hBD;
	13'h25C: q=8'hE7;
	13'h25D: q=8'hBE;
	13'h25E: q=8'hA6;
	13'h25F: q=8'h1;
	13'h260: q=8'hBD;
	13'h261: q=8'hE7;
	13'h262: q=8'hBE;
	13'h263: q=8'hCE;
	13'h264: q=8'hE1;
	13'h265: q=8'hAF;
	13'h266: q=8'hBD;
	13'h267: q=8'hE7;
	13'h268: q=8'hA8;
	13'h269: q=8'hDE;
	13'h26A: q=8'hE2;
	13'h26B: q=8'h8;
	13'h26C: q=8'h27;
	13'h26D: q=8'h3;
	13'h26E: q=8'hBD;
	13'h26F: q=8'hF4;
	13'h270: q=8'h12;
	13'h271: q=8'hBD;
	13'h272: q=8'hE7;
	13'h273: q=8'h6A;
	13'h274: q=8'hCE;
	13'h275: q=8'hE1;
	13'h276: q=8'hBC;
	13'h277: q=8'hBD;
	13'h278: q=8'hE7;
	13'h279: q=8'hA8;
	13'h27A: q=8'hCE;
	13'h27B: q=8'hFF;
	13'h27C: q=8'hFF;
	13'h27D: q=8'hDF;
	13'h27E: q=8'hE2;
	13'h27F: q=8'hBD;
	13'h280: q=8'hFA;
	13'h281: q=8'hA4;
	13'h282: q=8'h25;
	13'h283: q=8'hF6;
	13'h284: q=8'hDF;
	13'h285: q=8'hF4;
	13'h286: q=8'hBD;
	13'h287: q=8'h0;
	13'h288: q=8'hEB;
	13'h289: q=8'h27;
	13'h28A: q=8'hEF;
	13'h28B: q=8'h25;
	13'h28C: q=8'h6;
	13'h28D: q=8'hBD;
	13'h28E: q=8'hE3;
	13'h28F: q=8'h11;
	13'h290: q=8'h7E;
	13'h291: q=8'hE5;
	13'h292: q=8'h3D;
	13'h293: q=8'hBD;
	13'h294: q=8'hE6;
	13'h295: q=8'hB2;
	13'h296: q=8'hDE;
	13'h297: q=8'hA5;
	13'h298: q=8'hFF;
	13'h299: q=8'h42;
	13'h29A: q=8'hB0;
	13'h29B: q=8'hBD;
	13'h29C: q=8'hE3;
	13'h29D: q=8'h11;
	13'h29E: q=8'hD7;
	13'h29F: q=8'h82;
	13'h2A0: q=8'hBD;
	13'h2A1: q=8'hE3;
	13'h2A2: q=8'hB9;
	13'h2A3: q=8'h25;
	13'h2A4: q=8'h1C;
	13'h2A5: q=8'hDC;
	13'h2A6: q=8'hC1;
	13'h2A7: q=8'hA3;
	13'h2A8: q=8'h0;
	13'h2A9: q=8'hD3;
	13'h2AA: q=8'h95;
	13'h2AB: q=8'hDD;
	13'h2AC: q=8'h95;
	13'h2AD: q=8'h7;
	13'h2AE: q=8'h36;
	13'h2AF: q=8'h9F;
	13'h2B0: q=8'h91;
	13'h2B1: q=8'hF;
	13'h2B2: q=8'hAE;
	13'h2B3: q=8'h0;
	13'h2B4: q=8'h34;
	13'h2B5: q=8'h32;
	13'h2B6: q=8'hA7;
	13'h2B7: q=8'h0;
	13'h2B8: q=8'h8;
	13'h2B9: q=8'h9C;
	13'h2BA: q=8'h95;
	13'h2BB: q=8'h26;
	13'h2BC: q=8'hF8;
	13'h2BD: q=8'h9E;
	13'h2BE: q=8'h91;
	13'h2BF: q=8'h32;
	13'h2C0: q=8'h6;
	13'h2C1: q=8'hB6;
	13'h2C2: q=8'h42;
	13'h2C3: q=8'hB2;
	13'h2C4: q=8'h27;
	13'h2C5: q=8'h25;
	13'h2C6: q=8'hDC;
	13'h2C7: q=8'h95;
	13'h2C8: q=8'hDD;
	13'h2C9: q=8'hBD;
	13'h2CA: q=8'hDB;
	13'h2CB: q=8'h82;
	13'h2CC: q=8'h89;
	13'h2CD: q=8'h0;
	13'h2CE: q=8'hDD;
	13'h2CF: q=8'hBB;
	13'h2D0: q=8'hBD;
	13'h2D1: q=8'hE1;
	13'h2D2: q=8'hFE;
	13'h2D3: q=8'h7;
	13'h2D4: q=8'h36;
	13'h2D5: q=8'h9F;
	13'h2D6: q=8'h91;
	13'h2D7: q=8'hF;
	13'h2D8: q=8'h8E;
	13'h2D9: q=8'h42;
	13'h2DA: q=8'hAD;
	13'h2DB: q=8'h32;
	13'h2DC: q=8'hA7;
	13'h2DD: q=8'h0;
	13'h2DE: q=8'h8;
	13'h2DF: q=8'h9C;
	13'h2E0: q=8'hBF;
	13'h2E1: q=8'h26;
	13'h2E2: q=8'hF8;
	13'h2E3: q=8'h9E;
	13'h2E4: q=8'h91;
	13'h2E5: q=8'h32;
	13'h2E6: q=8'h6;
	13'h2E7: q=8'hDE;
	13'h2E8: q=8'hBB;
	13'h2E9: q=8'hDF;
	13'h2EA: q=8'h95;
	13'h2EB: q=8'hBD;
	13'h2EC: q=8'hE3;
	13'h2ED: q=8'hD9;
	13'h2EE: q=8'h8D;
	13'h2EF: q=8'h3;
	13'h2F0: q=8'h7E;
	13'h2F1: q=8'hE2;
	13'h2F2: q=8'h7A;
	13'h2F3: q=8'hDE;
	13'h2F4: q=8'h93;
	13'h2F5: q=8'hEC;
	13'h2F6: q=8'h0;
	13'h2F7: q=8'h26;
	13'h2F8: q=8'h1;
	13'h2F9: q=8'h39;
	13'h2FA: q=8'h3C;
	13'h2FB: q=8'hC6;
	13'h2FC: q=8'h4;
	13'h2FD: q=8'h3A;
	13'h2FE: q=8'h8;
	13'h2FF: q=8'hA6;
	13'h300: q=8'h0;
	13'h301: q=8'h26;
	13'h302: q=8'hFB;
	13'h303: q=8'h8;
	13'h304: q=8'h3C;
	13'h305: q=8'h30;
	13'h306: q=8'hEC;
	13'h307: q=8'h0;
	13'h308: q=8'hEE;
	13'h309: q=8'h2;
	13'h30A: q=8'hED;
	13'h30B: q=8'h0;
	13'h30C: q=8'h38;
	13'h30D: q=8'h31;
	13'h30E: q=8'h31;
	13'h30F: q=8'h20;
	13'h310: q=8'hE4;
	13'h311: q=8'h7F;
	13'h312: q=8'h0;
	13'h313: q=8'h85;
	13'h314: q=8'hDE;
	13'h315: q=8'hF4;
	13'h316: q=8'h9;
	13'h317: q=8'hDF;
	13'h318: q=8'hF4;
	13'h319: q=8'hCE;
	13'h31A: q=8'h42;
	13'h31B: q=8'hB1;
	13'h31C: q=8'hDF;
	13'h31D: q=8'hDE;
	13'h31E: q=8'h9F;
	13'h31F: q=8'h91;
	13'h320: q=8'h7;
	13'h321: q=8'h97;
	13'h322: q=8'h87;
	13'h323: q=8'h1;
	13'h324: q=8'hF;
	13'h325: q=8'h9E;
	13'h326: q=8'hF4;
	13'h327: q=8'h33;
	13'h328: q=8'hC1;
	13'h329: q=8'h20;
	13'h32A: q=8'h27;
	13'h32B: q=8'h38;
	13'h32C: q=8'hD7;
	13'h32D: q=8'h81;
	13'h32E: q=8'hC1;
	13'h32F: q=8'h22;
	13'h330: q=8'h27;
	13'h331: q=8'h5B;
	13'h332: q=8'h96;
	13'h333: q=8'h85;
	13'h334: q=8'h26;
	13'h335: q=8'h2E;
	13'h336: q=8'hC1;
	13'h337: q=8'h3F;
	13'h338: q=8'h26;
	13'h339: q=8'h4;
	13'h33A: q=8'hC6;
	13'h33B: q=8'h86;
	13'h33C: q=8'h20;
	13'h33D: q=8'h26;
	13'h33E: q=8'hC1;
	13'h33F: q=8'h30;
	13'h340: q=8'h25;
	13'h341: q=8'h4;
	13'h342: q=8'hC1;
	13'h343: q=8'h3C;
	13'h344: q=8'h25;
	13'h345: q=8'h1E;
	13'h346: q=8'h5D;
	13'h347: q=8'h2B;
	13'h348: q=8'h19;
	13'h349: q=8'hCE;
	13'h34A: q=8'hE0;
	13'h34B: q=8'h44;
	13'h34C: q=8'h9E;
	13'h34D: q=8'hF4;
	13'h34E: q=8'h5F;
	13'h34F: q=8'h8;
	13'h350: q=8'h32;
	13'h351: q=8'h81;
	13'h352: q=8'h20;
	13'h353: q=8'h27;
	13'h354: q=8'hFB;
	13'h355: q=8'hA0;
	13'h356: q=8'h0;
	13'h357: q=8'h27;
	13'h358: q=8'hF6;
	13'h359: q=8'h81;
	13'h35A: q=8'h80;
	13'h35B: q=8'h26;
	13'h35C: q=8'h35;
	13'h35D: q=8'hCA;
	13'h35E: q=8'h80;
	13'h35F: q=8'hDE;
	13'h360: q=8'hDE;
	13'h361: q=8'h8C;
	13'h362: q=8'hC6;
	13'h363: q=8'h21;
	13'h364: q=8'h9F;
	13'h365: q=8'hF4;
	13'h366: q=8'h9E;
	13'h367: q=8'h91;
	13'h368: q=8'h96;
	13'h369: q=8'h87;
	13'h36A: q=8'h6;
	13'h36B: q=8'h8;
	13'h36C: q=8'hDF;
	13'h36D: q=8'hDE;
	13'h36E: q=8'hE7;
	13'h36F: q=8'h0;
	13'h370: q=8'h27;
	13'h371: q=8'h38;
	13'h372: q=8'hC0;
	13'h373: q=8'h3A;
	13'h374: q=8'h27;
	13'h375: q=8'h4;
	13'h376: q=8'hC1;
	13'h377: q=8'h4B;
	13'h378: q=8'h26;
	13'h379: q=8'h2;
	13'h37A: q=8'hD7;
	13'h37B: q=8'h85;
	13'h37C: q=8'hC0;
	13'h37D: q=8'h49;
	13'h37E: q=8'h26;
	13'h37F: q=8'hA3;
	13'h380: q=8'hD7;
	13'h381: q=8'h81;
	13'h382: q=8'hF;
	13'h383: q=8'h9E;
	13'h384: q=8'hF4;
	13'h385: q=8'h33;
	13'h386: q=8'h5D;
	13'h387: q=8'h27;
	13'h388: q=8'hDB;
	13'h389: q=8'hD1;
	13'h38A: q=8'h81;
	13'h38B: q=8'h27;
	13'h38C: q=8'hD7;
	13'h38D: q=8'h8;
	13'h38E: q=8'hE7;
	13'h38F: q=8'h0;
	13'h390: q=8'h20;
	13'h391: q=8'hF3;
	13'h392: q=8'h9E;
	13'h393: q=8'hF4;
	13'h394: q=8'h5C;
	13'h395: q=8'hA6;
	13'h396: q=8'h0;
	13'h397: q=8'h8;
	13'h398: q=8'h2A;
	13'h399: q=8'hFB;
	13'h39A: q=8'hA6;
	13'h39B: q=8'h0;
	13'h39C: q=8'h26;
	13'h39D: q=8'hB2;
	13'h39E: q=8'h9F;
	13'h39F: q=8'hF4;
	13'h3A0: q=8'h9E;
	13'h3A1: q=8'h91;
	13'h3A2: q=8'hBD;
	13'h3A3: q=8'h42;
	13'h3A4: q=8'hA3;
	13'h3A5: q=8'h9E;
	13'h3A6: q=8'hF4;
	13'h3A7: q=8'h33;
	13'h3A8: q=8'h20;
	13'h3A9: q=8'hB5;
	13'h3AA: q=8'hE7;
	13'h3AB: q=8'h1;
	13'h3AC: q=8'hE7;
	13'h3AD: q=8'h2;
	13'h3AE: q=8'hDC;
	13'h3AF: q=8'hDE;
	13'h3B0: q=8'h83;
	13'h3B1: q=8'h42;
	13'h3B2: q=8'hAD;
	13'h3B3: q=8'hCE;
	13'h3B4: q=8'h42;
	13'h3B5: q=8'hB1;
	13'h3B6: q=8'hDF;
	13'h3B7: q=8'hF4;
	13'h3B8: q=8'h39;
	13'h3B9: q=8'hDE;
	13'h3BA: q=8'h93;
	13'h3BB: q=8'hEC;
	13'h3BC: q=8'h0;
	13'h3BD: q=8'h27;
	13'h3BE: q=8'hA;
	13'h3BF: q=8'hDC;
	13'h3C0: q=8'hA5;
	13'h3C1: q=8'hA3;
	13'h3C2: q=8'h2;
	13'h3C3: q=8'h23;
	13'h3C4: q=8'h5;
	13'h3C5: q=8'hEE;
	13'h3C6: q=8'h0;
	13'h3C7: q=8'h20;
	13'h3C8: q=8'hF2;
	13'h3C9: q=8'hD;
	13'h3CA: q=8'hDF;
	13'h3CB: q=8'hC1;
	13'h3CC: q=8'h39;
	13'h3CD: q=8'h26;
	13'h3CE: q=8'hFB;
	13'h3CF: q=8'hDE;
	13'h3D0: q=8'h93;
	13'h3D1: q=8'h6F;
	13'h3D2: q=8'h0;
	13'h3D3: q=8'h8;
	13'h3D4: q=8'h6F;
	13'h3D5: q=8'h0;
	13'h3D6: q=8'h8;
	13'h3D7: q=8'hDF;
	13'h3D8: q=8'h95;
	13'h3D9: q=8'hDE;
	13'h3DA: q=8'h93;
	13'h3DB: q=8'h9;
	13'h3DC: q=8'hDF;
	13'h3DD: q=8'hF4;
	13'h3DE: q=8'hBD;
	13'h3DF: q=8'h42;
	13'h3E0: q=8'h8E;
	13'h3E1: q=8'hDE;
	13'h3E2: q=8'hA1;
	13'h3E3: q=8'hDF;
	13'h3E4: q=8'h9D;
	13'h3E5: q=8'hBD;
	13'h3E6: q=8'hE5;
	13'h3E7: q=8'h60;
	13'h3E8: q=8'hDE;
	13'h3E9: q=8'h95;
	13'h3EA: q=8'hDF;
	13'h3EB: q=8'h97;
	13'h3EC: q=8'hDF;
	13'h3ED: q=8'h99;
	13'h3EE: q=8'hCE;
	13'h3EF: q=8'h42;
	13'h3F0: q=8'h41;
	13'h3F1: q=8'hFF;
	13'h3F2: q=8'h42;
	13'h3F3: q=8'h3D;
	13'h3F4: q=8'h38;
	13'h3F5: q=8'h9E;
	13'h3F6: q=8'h9B;
	13'h3F7: q=8'h4F;
	13'h3F8: q=8'h36;
	13'h3F9: q=8'h97;
	13'h3FA: q=8'hA7;
	13'h3FB: q=8'h97;
	13'h3FC: q=8'hA8;
	13'h3FD: q=8'h97;
	13'h3FE: q=8'h86;
	13'h3FF: q=8'hB7;
	13'h400: q=8'h42;
	13'h401: q=8'h6E;
	13'h402: q=8'h6E;
	13'h403: q=8'h0;
	13'h404: q=8'hC6;
	13'h405: q=8'hFE;
	13'h406: q=8'hD7;
	13'h407: q=8'hE8;
	13'h408: q=8'h7E;
	13'h409: q=8'h0;
	13'h40A: q=8'hF3;
	13'h40B: q=8'h8D;
	13'h40C: q=8'hF7;
	13'h40D: q=8'h7;
	13'h40E: q=8'h36;
	13'h40F: q=8'h8D;
	13'h410: q=8'hF7;
	13'h411: q=8'hBD;
	13'h412: q=8'hE6;
	13'h413: q=8'hB2;
	13'h414: q=8'h8D;
	13'h415: q=8'hA3;
	13'h416: q=8'h32;
	13'h417: q=8'h6;
	13'h418: q=8'h3C;
	13'h419: q=8'h27;
	13'h41A: q=8'h16;
	13'h41B: q=8'hBD;
	13'h41C: q=8'h0;
	13'h41D: q=8'hF3;
	13'h41E: q=8'h27;
	13'h41F: q=8'h16;
	13'h420: q=8'h81;
	13'h421: q=8'hA8;
	13'h422: q=8'h26;
	13'h423: q=8'hA;
	13'h424: q=8'hBD;
	13'h425: q=8'h0;
	13'h426: q=8'hEB;
	13'h427: q=8'h27;
	13'h428: q=8'h8;
	13'h429: q=8'hBD;
	13'h42A: q=8'hE6;
	13'h42B: q=8'hB2;
	13'h42C: q=8'h27;
	13'h42D: q=8'h8;
	13'h42E: q=8'h7E;
	13'h42F: q=8'hEA;
	13'h430: q=8'h3C;
	13'h431: q=8'hCE;
	13'h432: q=8'hFF;
	13'h433: q=8'hFF;
	13'h434: q=8'hDF;
	13'h435: q=8'hA5;
	13'h436: q=8'h38;
	13'h437: q=8'h31;
	13'h438: q=8'h31;
	13'h439: q=8'hBD;
	13'h43A: q=8'hE7;
	13'h43B: q=8'h6A;
	13'h43C: q=8'hBD;
	13'h43D: q=8'hE5;
	13'h43E: q=8'h66;
	13'h43F: q=8'hEC;
	13'h440: q=8'h0;
	13'h441: q=8'h26;
	13'h442: q=8'h6;
	13'h443: q=8'h7F;
	13'h444: q=8'h0;
	13'h445: q=8'hE8;
	13'h446: q=8'h7E;
	13'h447: q=8'hE2;
	13'h448: q=8'h71;
	13'h449: q=8'hEC;
	13'h44A: q=8'h2;
	13'h44B: q=8'h93;
	13'h44C: q=8'hA5;
	13'h44D: q=8'h22;
	13'h44E: q=8'hF4;
	13'h44F: q=8'hEC;
	13'h450: q=8'h2;
	13'h451: q=8'h3C;
	13'h452: q=8'hBD;
	13'h453: q=8'hF4;
	13'h454: q=8'h19;
	13'h455: q=8'h38;
	13'h456: q=8'h8;
	13'h457: q=8'h8;
	13'h458: q=8'h8;
	13'h459: q=8'h8;
	13'h45A: q=8'hDF;
	13'h45B: q=8'h89;
	13'h45C: q=8'h7F;
	13'h45D: q=8'h42;
	13'h45E: q=8'h84;
	13'h45F: q=8'h86;
	13'h460: q=8'h20;
	13'h461: q=8'h8C;
	13'h462: q=8'h86;
	13'h463: q=8'h21;
	13'h464: q=8'hDE;
	13'h465: q=8'h89;
	13'h466: q=8'h84;
	13'h467: q=8'h7F;
	13'h468: q=8'hBD;
	13'h469: q=8'hE7;
	13'h46A: q=8'hBE;
	13'h46B: q=8'hA6;
	13'h46C: q=8'h0;
	13'h46D: q=8'h8;
	13'h46E: q=8'h4D;
	13'h46F: q=8'h27;
	13'h470: q=8'hC8;
	13'h471: q=8'hF6;
	13'h472: q=8'h42;
	13'h473: q=8'h84;
	13'h474: q=8'h81;
	13'h475: q=8'h22;
	13'h476: q=8'h26;
	13'h477: q=8'h5;
	13'h478: q=8'hC8;
	13'h479: q=8'h1;
	13'h47A: q=8'hF7;
	13'h47B: q=8'h42;
	13'h47C: q=8'h84;
	13'h47D: q=8'h81;
	13'h47E: q=8'h3A;
	13'h47F: q=8'h26;
	13'h480: q=8'h9;
	13'h481: q=8'hC5;
	13'h482: q=8'h1;
	13'h483: q=8'h26;
	13'h484: q=8'h5;
	13'h485: q=8'hC4;
	13'h486: q=8'hFD;
	13'h487: q=8'hF7;
	13'h488: q=8'h42;
	13'h489: q=8'h84;
	13'h48A: q=8'h4D;
	13'h48B: q=8'h2A;
	13'h48C: q=8'hDB;
	13'h48D: q=8'h5D;
	13'h48E: q=8'h26;
	13'h48F: q=8'hD8;
	13'h490: q=8'h81;
	13'h491: q=8'h85;
	13'h492: q=8'h26;
	13'h493: q=8'h2;
	13'h494: q=8'hCA;
	13'h495: q=8'h2;
	13'h496: q=8'h81;
	13'h497: q=8'h83;
	13'h498: q=8'h26;
	13'h499: q=8'h2;
	13'h49A: q=8'hCA;
	13'h49B: q=8'h4;
	13'h49C: q=8'hF7;
	13'h49D: q=8'h42;
	13'h49E: q=8'h84;
	13'h49F: q=8'hBD;
	13'h4A0: q=8'h42;
	13'h4A1: q=8'hA6;
	13'h4A2: q=8'h81;
	13'h4A3: q=8'hC8;
	13'h4A4: q=8'h22;
	13'h4A5: q=8'hBC;
	13'h4A6: q=8'h8D;
	13'h4A7: q=8'hA;
	13'h4A8: q=8'hA6;
	13'h4A9: q=8'h0;
	13'h4AA: q=8'h2B;
	13'h4AB: q=8'hB8;
	13'h4AC: q=8'h8;
	13'h4AD: q=8'hBD;
	13'h4AE: q=8'hE7;
	13'h4AF: q=8'hBE;
	13'h4B0: q=8'h20;
	13'h4B1: q=8'hF6;
	13'h4B2: q=8'h80;
	13'h4B3: q=8'h7F;
	13'h4B4: q=8'hDF;
	13'h4B5: q=8'h89;
	13'h4B6: q=8'hCE;
	13'h4B7: q=8'hE0;
	13'h4B8: q=8'h45;
	13'h4B9: q=8'h4A;
	13'h4BA: q=8'h26;
	13'h4BB: q=8'h1;
	13'h4BC: q=8'h39;
	13'h4BD: q=8'h6D;
	13'h4BE: q=8'h0;
	13'h4BF: q=8'h8;
	13'h4C0: q=8'h2A;
	13'h4C1: q=8'hFB;
	13'h4C2: q=8'h20;
	13'h4C3: q=8'hF5;
	13'h4C4: q=8'h86;
	13'h4C5: q=8'h80;
	13'h4C6: q=8'h97;
	13'h4C7: q=8'h86;
	13'h4C8: q=8'hBD;
	13'h4C9: q=8'hE6;
	13'h4CA: q=8'hD3;
	13'h4CB: q=8'hBD;
	13'h4CC: q=8'hE1;
	13'h4CD: q=8'hD8;
	13'h4CE: q=8'h38;
	13'h4CF: q=8'h26;
	13'h4D0: q=8'h4;
	13'h4D1: q=8'hDE;
	13'h4D2: q=8'h89;
	13'h4D3: q=8'h3A;
	13'h4D4: q=8'h35;
	13'h4D5: q=8'hC6;
	13'h4D6: q=8'h9;
	13'h4D7: q=8'hBD;
	13'h4D8: q=8'hE2;
	13'h4D9: q=8'h1A;
	13'h4DA: q=8'hBD;
	13'h4DB: q=8'hE6;
	13'h4DC: q=8'h56;
	13'h4DD: q=8'h3C;
	13'h4DE: q=8'hDE;
	13'h4DF: q=8'hE2;
	13'h4E0: q=8'h3C;
	13'h4E1: q=8'hC6;
	13'h4E2: q=8'hA2;
	13'h4E3: q=8'hBD;
	13'h4E4: q=8'hEA;
	13'h4E5: q=8'h31;
	13'h4E6: q=8'hBD;
	13'h4E7: q=8'hE9;
	13'h4E8: q=8'hE;
	13'h4E9: q=8'hBD;
	13'h4EA: q=8'hE9;
	13'h4EB: q=8'hC;
	13'h4EC: q=8'hD6;
	13'h4ED: q=8'hCE;
	13'h4EE: q=8'hCA;
	13'h4EF: q=8'h7F;
	13'h4F0: q=8'hD4;
	13'h4F1: q=8'hCA;
	13'h4F2: q=8'hD7;
	13'h4F3: q=8'hCA;
	13'h4F4: q=8'hCE;
	13'h4F5: q=8'hE4;
	13'h4F6: q=8'hFA;
	13'h4F7: q=8'h7E;
	13'h4F8: q=8'hE9;
	13'h4F9: q=8'hA4;
	13'h4FA: q=8'hCE;
	13'h4FB: q=8'hF0;
	13'h4FC: q=8'h8B;
	13'h4FD: q=8'hBD;
	13'h4FE: q=8'hF2;
	13'h4FF: q=8'h51;
	13'h500: q=8'hBD;
	13'h501: q=8'h0;
	13'h502: q=8'hF3;
	13'h503: q=8'h81;
	13'h504: q=8'hA5;
	13'h505: q=8'h26;
	13'h506: q=8'h6;
	13'h507: q=8'hBD;
	13'h508: q=8'h0;
	13'h509: q=8'hEB;
	13'h50A: q=8'hBD;
	13'h50B: q=8'hE9;
	13'h50C: q=8'hC;
	13'h50D: q=8'hBD;
	13'h50E: q=8'hF2;
	13'h50F: q=8'hAD;
	13'h510: q=8'hBD;
	13'h511: q=8'hE9;
	13'h512: q=8'hA2;
	13'h513: q=8'hDE;
	13'h514: q=8'hB5;
	13'h515: q=8'h3C;
	13'h516: q=8'h86;
	13'h517: q=8'h80;
	13'h518: q=8'h36;
	13'h519: q=8'h8D;
	13'h51A: q=8'h4B;
	13'h51B: q=8'hDE;
	13'h51C: q=8'hF4;
	13'h51D: q=8'hDF;
	13'h51E: q=8'hA9;
	13'h51F: q=8'hA6;
	13'h520: q=8'h0;
	13'h521: q=8'h27;
	13'h522: q=8'h7;
	13'h523: q=8'h81;
	13'h524: q=8'h3A;
	13'h525: q=8'h27;
	13'h526: q=8'h16;
	13'h527: q=8'h7E;
	13'h528: q=8'hEA;
	13'h529: q=8'h3C;
	13'h52A: q=8'h8;
	13'h52B: q=8'hA6;
	13'h52C: q=8'h0;
	13'h52D: q=8'h8;
	13'h52E: q=8'hAA;
	13'h52F: q=8'h0;
	13'h530: q=8'hB7;
	13'h531: q=8'h42;
	13'h532: q=8'h83;
	13'h533: q=8'h27;
	13'h534: q=8'h54;
	13'h535: q=8'h8;
	13'h536: q=8'hEC;
	13'h537: q=8'h0;
	13'h538: q=8'hDD;
	13'h539: q=8'hE2;
	13'h53A: q=8'h8;
	13'h53B: q=8'hDF;
	13'h53C: q=8'hF4;
	13'h53D: q=8'hBD;
	13'h53E: q=8'h0;
	13'h53F: q=8'hEB;
	13'h540: q=8'h8D;
	13'h541: q=8'h2;
	13'h542: q=8'h20;
	13'h543: q=8'hD5;
	13'h544: q=8'h27;
	13'h545: q=8'h71;
	13'h546: q=8'hBD;
	13'h547: q=8'h42;
	13'h548: q=8'hA0;
	13'h549: q=8'h4D;
	13'h54A: q=8'h2B;
	13'h54B: q=8'h3;
	13'h54C: q=8'h7E;
	13'h54D: q=8'hE6;
	13'h54E: q=8'hD3;
	13'h54F: q=8'h81;
	13'h550: q=8'hA0;
	13'h551: q=8'h22;
	13'h552: q=8'hD4;
	13'h553: q=8'h48;
	13'h554: q=8'h16;
	13'h555: q=8'hCE;
	13'h556: q=8'hE1;
	13'h557: q=8'h48;
	13'h558: q=8'h3A;
	13'h559: q=8'hEE;
	13'h55A: q=8'h0;
	13'h55B: q=8'hBD;
	13'h55C: q=8'h0;
	13'h55D: q=8'hEB;
	13'h55E: q=8'h6E;
	13'h55F: q=8'h0;
	13'h560: q=8'hDE;
	13'h561: q=8'h93;
	13'h562: q=8'h9;
	13'h563: q=8'hDF;
	13'h564: q=8'hAD;
	13'h565: q=8'h39;
	13'h566: q=8'hBD;
	13'h567: q=8'hF8;
	13'h568: q=8'h79;
	13'h569: q=8'h27;
	13'h56A: q=8'hB;
	13'h56B: q=8'h81;
	13'h56C: q=8'h3;
	13'h56D: q=8'h27;
	13'h56E: q=8'hF;
	13'h56F: q=8'h81;
	13'h570: q=8'h13;
	13'h571: q=8'h27;
	13'h572: q=8'h4;
	13'h573: q=8'hB7;
	13'h574: q=8'h42;
	13'h575: q=8'h7F;
	13'h576: q=8'h39;
	13'h577: q=8'hBD;
	13'h578: q=8'hF8;
	13'h579: q=8'h83;
	13'h57A: q=8'h27;
	13'h57B: q=8'hFB;
	13'h57C: q=8'h20;
	13'h57D: q=8'hED;
	13'h57E: q=8'hD;
	13'h57F: q=8'h26;
	13'h580: q=8'h36;
	13'h581: q=8'hDE;
	13'h582: q=8'hF4;
	13'h583: q=8'hDF;
	13'h584: q=8'hA9;
	13'h585: q=8'h76;
	13'h586: q=8'h42;
	13'h587: q=8'h83;
	13'h588: q=8'h38;
	13'h589: q=8'hDE;
	13'h58A: q=8'hE2;
	13'h58B: q=8'h8;
	13'h58C: q=8'h27;
	13'h58D: q=8'h7;
	13'h58E: q=8'h9;
	13'h58F: q=8'hDF;
	13'h590: q=8'hA3;
	13'h591: q=8'hDE;
	13'h592: q=8'hA9;
	13'h593: q=8'hDF;
	13'h594: q=8'hA7;
	13'h595: q=8'h7F;
	13'h596: q=8'h0;
	13'h597: q=8'hE8;
	13'h598: q=8'hCE;
	13'h599: q=8'hE1;
	13'h59A: q=8'hC0;
	13'h59B: q=8'h7D;
	13'h59C: q=8'h42;
	13'h59D: q=8'h83;
	13'h59E: q=8'h2A;
	13'h59F: q=8'h3;
	13'h5A0: q=8'h7E;
	13'h5A1: q=8'hE2;
	13'h5A2: q=8'h66;
	13'h5A3: q=8'h7E;
	13'h5A4: q=8'hE2;
	13'h5A5: q=8'h71;
	13'h5A6: q=8'h26;
	13'h5A7: q=8'hF;
	13'h5A8: q=8'hC6;
	13'h5A9: q=8'h20;
	13'h5AA: q=8'hDE;
	13'h5AB: q=8'hA7;
	13'h5AC: q=8'h26;
	13'h5AD: q=8'h3;
	13'h5AE: q=8'h7E;
	13'h5AF: q=8'hE2;
	13'h5B0: q=8'h38;
	13'h5B1: q=8'hDF;
	13'h5B2: q=8'hF4;
	13'h5B3: q=8'hDE;
	13'h5B4: q=8'hA3;
	13'h5B5: q=8'hDF;
	13'h5B6: q=8'hE2;
	13'h5B7: q=8'h39;
	13'h5B8: q=8'h27;
	13'h5B9: q=8'h3A;
	13'h5BA: q=8'hBD;
	13'h5BB: q=8'hEB;
	13'h5BC: q=8'hBD;
	13'h5BD: q=8'h37;
	13'h5BE: q=8'h36;
	13'h5BF: q=8'hDE;
	13'h5C0: q=8'hA1;
	13'h5C1: q=8'hDF;
	13'h5C2: q=8'hCC;
	13'h5C3: q=8'hBD;
	13'h5C4: q=8'h0;
	13'h5C5: q=8'hF3;
	13'h5C6: q=8'h27;
	13'h5C7: q=8'h12;
	13'h5C8: q=8'hBD;
	13'h5C9: q=8'hEA;
	13'h5CA: q=8'h2F;
	13'h5CB: q=8'hBD;
	13'h5CC: q=8'hEF;
	13'h5CD: q=8'h4C;
	13'h5CE: q=8'hDE;
	13'h5CF: q=8'hCC;
	13'h5D0: q=8'h9;
	13'h5D1: q=8'hDF;
	13'h5D2: q=8'hCC;
	13'h5D3: q=8'hFC;
	13'h5D4: q=8'h42;
	13'h5D5: q=8'h50;
	13'h5D6: q=8'h93;
	13'h5D7: q=8'hCC;
	13'h5D8: q=8'h25;
	13'h5D9: q=8'h1D;
	13'h5DA: q=8'hDC;
	13'h5DB: q=8'hCC;
	13'h5DC: q=8'h37;
	13'h5DD: q=8'h36;
	13'h5DE: q=8'h30;
	13'h5DF: q=8'hA3;
	13'h5E0: q=8'h2;
	13'h5E1: q=8'h25;
	13'h5E2: q=8'h14;
	13'h5E3: q=8'hED;
	13'h5E4: q=8'h2;
	13'h5E5: q=8'h83;
	13'h5E6: q=8'h0;
	13'h5E7: q=8'h3A;
	13'h5E8: q=8'h25;
	13'h5E9: q=8'hD;
	13'h5EA: q=8'h93;
	13'h5EB: q=8'h95;
	13'h5EC: q=8'h25;
	13'h5ED: q=8'h9;
	13'h5EE: q=8'h38;
	13'h5EF: q=8'hDF;
	13'h5F0: q=8'hA1;
	13'h5F1: q=8'h38;
	13'h5F2: q=8'hDF;
	13'h5F3: q=8'h9B;
	13'h5F4: q=8'h7E;
	13'h5F5: q=8'hE3;
	13'h5F6: q=8'hDE;
	13'h5F7: q=8'h7E;
	13'h5F8: q=8'hE2;
	13'h5F9: q=8'h36;
	13'h5FA: q=8'h26;
	13'h5FB: q=8'h3;
	13'h5FC: q=8'h7E;
	13'h5FD: q=8'hE3;
	13'h5FE: q=8'hD9;
	13'h5FF: q=8'hBD;
	13'h600: q=8'hE3;
	13'h601: q=8'hDE;
	13'h602: q=8'h20;
	13'h603: q=8'hE;
	13'h604: q=8'hC6;
	13'h605: q=8'h3;
	13'h606: q=8'hBD;
	13'h607: q=8'hE2;
	13'h608: q=8'h1A;
	13'h609: q=8'hDE;
	13'h60A: q=8'hF4;
	13'h60B: q=8'h3C;
	13'h60C: q=8'hDE;
	13'h60D: q=8'hE2;
	13'h60E: q=8'h3C;
	13'h60F: q=8'h86;
	13'h610: q=8'h82;
	13'h611: q=8'h36;
	13'h612: q=8'hBD;
	13'h613: q=8'h0;
	13'h614: q=8'hF3;
	13'h615: q=8'h8D;
	13'h616: q=8'h3;
	13'h617: q=8'h7E;
	13'h618: q=8'hE5;
	13'h619: q=8'h19;
	13'h61A: q=8'hBD;
	13'h61B: q=8'hE6;
	13'h61C: q=8'hB2;
	13'h61D: q=8'h8D;
	13'h61E: q=8'h3A;
	13'h61F: q=8'h8;
	13'h620: q=8'hDC;
	13'h621: q=8'hA5;
	13'h622: q=8'h93;
	13'h623: q=8'hE2;
	13'h624: q=8'h22;
	13'h625: q=8'h2;
	13'h626: q=8'hDE;
	13'h627: q=8'h93;
	13'h628: q=8'hBD;
	13'h629: q=8'hE3;
	13'h62A: q=8'hBB;
	13'h62B: q=8'h25;
	13'h62C: q=8'h15;
	13'h62D: q=8'h9;
	13'h62E: q=8'hDF;
	13'h62F: q=8'hF4;
	13'h630: q=8'h39;
	13'h631: q=8'h26;
	13'h632: q=8'hFD;
	13'h633: q=8'h86;
	13'h634: q=8'hFF;
	13'h635: q=8'h97;
	13'h636: q=8'hB5;
	13'h637: q=8'hBD;
	13'h638: q=8'hE1;
	13'h639: q=8'hD8;
	13'h63A: q=8'h35;
	13'h63B: q=8'h81;
	13'h63C: q=8'h2;
	13'h63D: q=8'h27;
	13'h63E: q=8'hB;
	13'h63F: q=8'hC6;
	13'h640: q=8'h4;
	13'h641: q=8'h8C;
	13'h642: q=8'hC6;
	13'h643: q=8'hE;
	13'h644: q=8'h7E;
	13'h645: q=8'hE2;
	13'h646: q=8'h38;
	13'h647: q=8'h7E;
	13'h648: q=8'hEA;
	13'h649: q=8'h3C;
	13'h64A: q=8'h32;
	13'h64B: q=8'h38;
	13'h64C: q=8'hDF;
	13'h64D: q=8'hE2;
	13'h64E: q=8'h38;
	13'h64F: q=8'hDF;
	13'h650: q=8'hF4;
	13'h651: q=8'h8D;
	13'h652: q=8'h3;
	13'h653: q=8'hDF;
	13'h654: q=8'hF4;
	13'h655: q=8'h39;
	13'h656: q=8'hC6;
	13'h657: q=8'h3A;
	13'h658: q=8'h86;
	13'h659: q=8'h5F;
	13'h65A: q=8'hD7;
	13'h65B: q=8'h80;
	13'h65C: q=8'h5F;
	13'h65D: q=8'hDE;
	13'h65E: q=8'hF4;
	13'h65F: q=8'h17;
	13'h660: q=8'hD6;
	13'h661: q=8'h80;
	13'h662: q=8'h97;
	13'h663: q=8'h80;
	13'h664: q=8'hA6;
	13'h665: q=8'h0;
	13'h666: q=8'h27;
	13'h667: q=8'hED;
	13'h668: q=8'h11;
	13'h669: q=8'h27;
	13'h66A: q=8'hEA;
	13'h66B: q=8'h8;
	13'h66C: q=8'h81;
	13'h66D: q=8'h22;
	13'h66E: q=8'h27;
	13'h66F: q=8'hEF;
	13'h670: q=8'h20;
	13'h671: q=8'hF2;
	13'h672: q=8'hBD;
	13'h673: q=8'hE9;
	13'h674: q=8'hC;
	13'h675: q=8'hBD;
	13'h676: q=8'h0;
	13'h677: q=8'hF3;
	13'h678: q=8'h81;
	13'h679: q=8'h81;
	13'h67A: q=8'h27;
	13'h67B: q=8'h5;
	13'h67C: q=8'hC6;
	13'h67D: q=8'hA3;
	13'h67E: q=8'hBD;
	13'h67F: q=8'hEA;
	13'h680: q=8'h31;
	13'h681: q=8'h96;
	13'h682: q=8'hC9;
	13'h683: q=8'h26;
	13'h684: q=8'h5;
	13'h685: q=8'h8D;
	13'h686: q=8'hD2;
	13'h687: q=8'hDF;
	13'h688: q=8'hF4;
	13'h689: q=8'h39;
	13'h68A: q=8'hBD;
	13'h68B: q=8'h0;
	13'h68C: q=8'hF3;
	13'h68D: q=8'h25;
	13'h68E: q=8'h8B;
	13'h68F: q=8'h7E;
	13'h690: q=8'hE5;
	13'h691: q=8'h44;
	13'h692: q=8'hBD;
	13'h693: q=8'hEF;
	13'h694: q=8'hD;
	13'h695: q=8'h36;
	13'h696: q=8'h81;
	13'h697: q=8'h82;
	13'h698: q=8'h27;
	13'h699: q=8'h4;
	13'h69A: q=8'h81;
	13'h69B: q=8'h81;
	13'h69C: q=8'h26;
	13'h69D: q=8'hA9;
	13'h69E: q=8'h7A;
	13'h69F: q=8'h0;
	13'h6A0: q=8'hCD;
	13'h6A1: q=8'h26;
	13'h6A2: q=8'h4;
	13'h6A3: q=8'h32;
	13'h6A4: q=8'h7E;
	13'h6A5: q=8'hE5;
	13'h6A6: q=8'h46;
	13'h6A7: q=8'hBD;
	13'h6A8: q=8'h0;
	13'h6A9: q=8'hEB;
	13'h6AA: q=8'h8D;
	13'h6AB: q=8'h6;
	13'h6AC: q=8'h81;
	13'h6AD: q=8'h2C;
	13'h6AE: q=8'h27;
	13'h6AF: q=8'hEE;
	13'h6B0: q=8'h31;
	13'h6B1: q=8'h39;
	13'h6B2: q=8'hCE;
	13'h6B3: q=8'h0;
	13'h6B4: q=8'h0;
	13'h6B5: q=8'hDF;
	13'h6B6: q=8'hA5;
	13'h6B7: q=8'h24;
	13'h6B8: q=8'hF8;
	13'h6B9: q=8'h80;
	13'h6BA: q=8'h30;
	13'h6BB: q=8'h97;
	13'h6BC: q=8'h80;
	13'h6BD: q=8'hDC;
	13'h6BE: q=8'hA5;
	13'h6BF: q=8'h81;
	13'h6C0: q=8'h18;
	13'h6C1: q=8'h22;
	13'h6C2: q=8'hD9;
	13'h6C3: q=8'h5;
	13'h6C4: q=8'h5;
	13'h6C5: q=8'hD3;
	13'h6C6: q=8'hA5;
	13'h6C7: q=8'h5;
	13'h6C8: q=8'hDB;
	13'h6C9: q=8'h80;
	13'h6CA: q=8'h89;
	13'h6CB: q=8'h0;
	13'h6CC: q=8'hDD;
	13'h6CD: q=8'hA5;
	13'h6CE: q=8'hBD;
	13'h6CF: q=8'h0;
	13'h6D0: q=8'hEB;
	13'h6D1: q=8'h20;
	13'h6D2: q=8'hE4;
	13'h6D3: q=8'hBD;
	13'h6D4: q=8'hEB;
	13'h6D5: q=8'h1B;
	13'h6D6: q=8'hDF;
	13'h6D7: q=8'hB5;
	13'h6D8: q=8'hC6;
	13'h6D9: q=8'hAF;
	13'h6DA: q=8'hBD;
	13'h6DB: q=8'hEA;
	13'h6DC: q=8'h31;
	13'h6DD: q=8'h96;
	13'h6DE: q=8'h84;
	13'h6DF: q=8'h36;
	13'h6E0: q=8'hBD;
	13'h6E1: q=8'hE9;
	13'h6E2: q=8'h1A;
	13'h6E3: q=8'h32;
	13'h6E4: q=8'h46;
	13'h6E5: q=8'hBD;
	13'h6E6: q=8'hE9;
	13'h6E7: q=8'h10;
	13'h6E8: q=8'h27;
	13'h6E9: q=8'h2F;
	13'h6EA: q=8'hDE;
	13'h6EB: q=8'hCC;
	13'h6EC: q=8'hDC;
	13'h6ED: q=8'h9B;
	13'h6EE: q=8'hA3;
	13'h6EF: q=8'h2;
	13'h6F0: q=8'h24;
	13'h6F1: q=8'h13;
	13'h6F2: q=8'hDC;
	13'h6F3: q=8'h95;
	13'h6F4: q=8'h93;
	13'h6F5: q=8'hCC;
	13'h6F6: q=8'h22;
	13'h6F7: q=8'hD;
	13'h6F8: q=8'hE6;
	13'h6F9: q=8'h0;
	13'h6FA: q=8'hBD;
	13'h6FB: q=8'hEC;
	13'h6FC: q=8'hFC;
	13'h6FD: q=8'hDE;
	13'h6FE: q=8'hC7;
	13'h6FF: q=8'hBD;
	13'h700: q=8'hEE;
	13'h701: q=8'h38;
	13'h702: q=8'hCE;
	13'h703: q=8'h0;
	13'h704: q=8'hD0;
	13'h705: q=8'hDF;
	13'h706: q=8'hC7;
	13'h707: q=8'hBD;
	13'h708: q=8'hEE;
	13'h709: q=8'h70;
	13'h70A: q=8'hDE;
	13'h70B: q=8'hC7;
	13'h70C: q=8'hA6;
	13'h70D: q=8'h0;
	13'h70E: q=8'h36;
	13'h70F: q=8'hEC;
	13'h710: q=8'h2;
	13'h711: q=8'hDE;
	13'h712: q=8'hB5;
	13'h713: q=8'hED;
	13'h714: q=8'h2;
	13'h715: q=8'h32;
	13'h716: q=8'hA7;
	13'h717: q=8'h0;
	13'h718: q=8'h39;
	13'h719: q=8'h7E;
	13'h71A: q=8'hF2;
	13'h71B: q=8'h70;
	13'h71C: q=8'hBD;
	13'h71D: q=8'hE4;
	13'h71E: q=8'h4;
	13'h71F: q=8'h8D;
	13'h720: q=8'h4;
	13'h721: q=8'h7F;
	13'h722: q=8'h0;
	13'h723: q=8'hE8;
	13'h724: q=8'h39;
	13'h725: q=8'h27;
	13'h726: q=8'h3F;
	13'h727: q=8'h81;
	13'h728: q=8'h40;
	13'h729: q=8'h26;
	13'h72A: q=8'hB;
	13'h72B: q=8'hBD;
	13'h72C: q=8'hFC;
	13'h72D: q=8'h29;
	13'h72E: q=8'hBD;
	13'h72F: q=8'h0;
	13'h730: q=8'hF3;
	13'h731: q=8'h27;
	13'h732: q=8'h33;
	13'h733: q=8'hBD;
	13'h734: q=8'hEA;
	13'h735: q=8'h2F;
	13'h736: q=8'h27;
	13'h737: q=8'h3B;
	13'h738: q=8'h81;
	13'h739: q=8'hA1;
	13'h73A: q=8'h27;
	13'h73B: q=8'h50;
	13'h73C: q=8'h81;
	13'h73D: q=8'h2C;
	13'h73E: q=8'h27;
	13'h73F: q=8'h34;
	13'h740: q=8'h81;
	13'h741: q=8'h3B;
	13'h742: q=8'h27;
	13'h743: q=8'h5E;
	13'h744: q=8'hBD;
	13'h745: q=8'hE9;
	13'h746: q=8'h1A;
	13'h747: q=8'h96;
	13'h748: q=8'h84;
	13'h749: q=8'h36;
	13'h74A: q=8'h26;
	13'h74B: q=8'h6;
	13'h74C: q=8'hBD;
	13'h74D: q=8'hF4;
	13'h74E: q=8'h26;
	13'h74F: q=8'hBD;
	13'h750: q=8'hED;
	13'h751: q=8'h5;
	13'h752: q=8'h8D;
	13'h753: q=8'h57;
	13'h754: q=8'h33;
	13'h755: q=8'h5D;
	13'h756: q=8'h26;
	13'h757: q=8'h9;
	13'h758: q=8'hBD;
	13'h759: q=8'h0;
	13'h75A: q=8'hF3;
	13'h75B: q=8'h81;
	13'h75C: q=8'h2C;
	13'h75D: q=8'h27;
	13'h75E: q=8'h15;
	13'h75F: q=8'h8D;
	13'h760: q=8'h58;
	13'h761: q=8'hBD;
	13'h762: q=8'h0;
	13'h763: q=8'hF3;
	13'h764: q=8'h26;
	13'h765: q=8'hD2;
	13'h766: q=8'h86;
	13'h767: q=8'hD;
	13'h768: q=8'h20;
	13'h769: q=8'h54;
	13'h76A: q=8'hBD;
	13'h76B: q=8'hFA;
	13'h76C: q=8'h7B;
	13'h76D: q=8'h27;
	13'h76E: q=8'hF7;
	13'h76F: q=8'h96;
	13'h770: q=8'hE6;
	13'h771: q=8'h26;
	13'h772: q=8'hF3;
	13'h773: q=8'h39;
	13'h774: q=8'hBD;
	13'h775: q=8'hFA;
	13'h776: q=8'h7B;
	13'h777: q=8'h27;
	13'h778: q=8'hA;
	13'h779: q=8'hD6;
	13'h77A: q=8'hE6;
	13'h77B: q=8'hD1;
	13'h77C: q=8'hE5;
	13'h77D: q=8'h25;
	13'h77E: q=8'h6;
	13'h77F: q=8'h8D;
	13'h780: q=8'hE5;
	13'h781: q=8'h20;
	13'h782: q=8'h1F;
	13'h783: q=8'hD6;
	13'h784: q=8'hE6;
	13'h785: q=8'hD0;
	13'h786: q=8'hE4;
	13'h787: q=8'h24;
	13'h788: q=8'hFC;
	13'h789: q=8'h50;
	13'h78A: q=8'h20;
	13'h78B: q=8'h11;
	13'h78C: q=8'hBD;
	13'h78D: q=8'hEF;
	13'h78E: q=8'hA;
	13'h78F: q=8'h81;
	13'h790: q=8'h29;
	13'h791: q=8'h27;
	13'h792: q=8'h3;
	13'h793: q=8'h7E;
	13'h794: q=8'hEA;
	13'h795: q=8'h3C;
	13'h796: q=8'hBD;
	13'h797: q=8'hFA;
	13'h798: q=8'h7B;
	13'h799: q=8'hD0;
	13'h79A: q=8'hE6;
	13'h79B: q=8'h23;
	13'h79C: q=8'h5;
	13'h79D: q=8'h8D;
	13'h79E: q=8'h1A;
	13'h79F: q=8'h5A;
	13'h7A0: q=8'h26;
	13'h7A1: q=8'hFB;
	13'h7A2: q=8'hBD;
	13'h7A3: q=8'h0;
	13'h7A4: q=8'hEB;
	13'h7A5: q=8'h7E;
	13'h7A6: q=8'hE7;
	13'h7A7: q=8'h36;
	13'h7A8: q=8'hBD;
	13'h7A9: q=8'hED;
	13'h7AA: q=8'h6;
	13'h7AB: q=8'hBD;
	13'h7AC: q=8'hEE;
	13'h7AD: q=8'h56;
	13'h7AE: q=8'h5C;
	13'h7AF: q=8'h5A;
	13'h7B0: q=8'h27;
	13'h7B1: q=8'hC1;
	13'h7B2: q=8'hA6;
	13'h7B3: q=8'h0;
	13'h7B4: q=8'h8;
	13'h7B5: q=8'h8D;
	13'h7B6: q=8'h7;
	13'h7B7: q=8'h20;
	13'h7B8: q=8'hF6;
	13'h7B9: q=8'h86;
	13'h7BA: q=8'h20;
	13'h7BB: q=8'h8C;
	13'h7BC: q=8'h86;
	13'h7BD: q=8'h3F;
	13'h7BE: q=8'h7E;
	13'h7BF: q=8'hF9;
	13'h7C0: q=8'hC6;
	13'h7C1: q=8'h3F;
	13'h7C2: q=8'h52;
	13'h7C3: q=8'h45;
	13'h7C4: q=8'h44;
	13'h7C5: q=8'h4F;
	13'h7C6: q=8'hD;
	13'h7C7: q=8'h0;
	13'h7C8: q=8'h96;
	13'h7C9: q=8'h87;
	13'h7CA: q=8'h27;
	13'h7CB: q=8'h7;
	13'h7CC: q=8'hDE;
	13'h7CD: q=8'hAB;
	13'h7CE: q=8'hDF;
	13'h7CF: q=8'hE2;
	13'h7D0: q=8'h7E;
	13'h7D1: q=8'hEA;
	13'h7D2: q=8'h3C;
	13'h7D3: q=8'hCE;
	13'h7D4: q=8'hE7;
	13'h7D5: q=8'hC0;
	13'h7D6: q=8'hBD;
	13'h7D7: q=8'hE7;
	13'h7D8: q=8'hA8;
	13'h7D9: q=8'hDE;
	13'h7DA: q=8'hA9;
	13'h7DB: q=8'hDF;
	13'h7DC: q=8'hF4;
	13'h7DD: q=8'h39;
	13'h7DE: q=8'hC6;
	13'h7DF: q=8'h16;
	13'h7E0: q=8'hDE;
	13'h7E1: q=8'hE2;
	13'h7E2: q=8'h8;
	13'h7E3: q=8'h26;
	13'h7E4: q=8'h3;
	13'h7E5: q=8'h7E;
	13'h7E6: q=8'hE2;
	13'h7E7: q=8'h38;
	13'h7E8: q=8'h81;
	13'h7E9: q=8'h22;
	13'h7EA: q=8'h26;
	13'h7EB: q=8'hB;
	13'h7EC: q=8'hBD;
	13'h7ED: q=8'hEA;
	13'h7EE: q=8'h7;
	13'h7EF: q=8'hC6;
	13'h7F0: q=8'h3B;
	13'h7F1: q=8'hBD;
	13'h7F2: q=8'hEA;
	13'h7F3: q=8'h31;
	13'h7F4: q=8'hBD;
	13'h7F5: q=8'hE7;
	13'h7F6: q=8'hAB;
	13'h7F7: q=8'h8D;
	13'h7F8: q=8'h6;
	13'h7F9: q=8'hC6;
	13'h7FA: q=8'h2C;
	13'h7FB: q=8'hE7;
	13'h7FC: q=8'h0;
	13'h7FD: q=8'h20;
	13'h7FE: q=8'h12;
	13'h7FF: q=8'hBD;
	13'h800: q=8'hE7;
	13'h801: q=8'hBC;
	13'h802: q=8'hBD;
	13'h803: q=8'hE7;
	13'h804: q=8'hB9;
	13'h805: q=8'hBD;
	13'h806: q=8'hFA;
	13'h807: q=8'hA4;
	13'h808: q=8'h24;
	13'h809: q=8'hD3;
	13'h80A: q=8'h38;
	13'h80B: q=8'h7E;
	13'h80C: q=8'hE5;
	13'h80D: q=8'h85;
	13'h80E: q=8'hDE;
	13'h80F: q=8'hAD;
	13'h810: q=8'h86;
	13'h811: q=8'h4F;
	13'h812: q=8'h97;
	13'h813: q=8'h87;
	13'h814: q=8'hDF;
	13'h815: q=8'hAF;
	13'h816: q=8'hBD;
	13'h817: q=8'hEB;
	13'h818: q=8'h1B;
	13'h819: q=8'hDF;
	13'h81A: q=8'hB5;
	13'h81B: q=8'hDE;
	13'h81C: q=8'hF4;
	13'h81D: q=8'hDF;
	13'h81E: q=8'hA5;
	13'h81F: q=8'hDE;
	13'h820: q=8'hAF;
	13'h821: q=8'hA6;
	13'h822: q=8'h0;
	13'h823: q=8'h26;
	13'h824: q=8'h9;
	13'h825: q=8'h96;
	13'h826: q=8'h87;
	13'h827: q=8'h26;
	13'h828: q=8'h4E;
	13'h829: q=8'hBD;
	13'h82A: q=8'hE7;
	13'h82B: q=8'hBC;
	13'h82C: q=8'h8D;
	13'h82D: q=8'hD1;
	13'h82E: q=8'hDF;
	13'h82F: q=8'hF4;
	13'h830: q=8'hBD;
	13'h831: q=8'h0;
	13'h832: q=8'hEB;
	13'h833: q=8'hD6;
	13'h834: q=8'h84;
	13'h835: q=8'h27;
	13'h836: q=8'h1C;
	13'h837: q=8'hDE;
	13'h838: q=8'hF4;
	13'h839: q=8'h97;
	13'h83A: q=8'h80;
	13'h83B: q=8'h81;
	13'h83C: q=8'h22;
	13'h83D: q=8'h27;
	13'h83E: q=8'h7;
	13'h83F: q=8'h9;
	13'h840: q=8'h86;
	13'h841: q=8'h3A;
	13'h842: q=8'h97;
	13'h843: q=8'h80;
	13'h844: q=8'h86;
	13'h845: q=8'h2C;
	13'h846: q=8'h97;
	13'h847: q=8'h81;
	13'h848: q=8'hBD;
	13'h849: q=8'hED;
	13'h84A: q=8'hC;
	13'h84B: q=8'hBD;
	13'h84C: q=8'hEF;
	13'h84D: q=8'h3E;
	13'h84E: q=8'hBD;
	13'h84F: q=8'hE6;
	13'h850: q=8'hEA;
	13'h851: q=8'h20;
	13'h852: q=8'h6;
	13'h853: q=8'hBD;
	13'h854: q=8'hF3;
	13'h855: q=8'h59;
	13'h856: q=8'hBD;
	13'h857: q=8'hF2;
	13'h858: q=8'h70;
	13'h859: q=8'hBD;
	13'h85A: q=8'h0;
	13'h85B: q=8'hF3;
	13'h85C: q=8'h27;
	13'h85D: q=8'h7;
	13'h85E: q=8'h81;
	13'h85F: q=8'h2C;
	13'h860: q=8'h27;
	13'h861: q=8'h3;
	13'h862: q=8'h7E;
	13'h863: q=8'hE7;
	13'h864: q=8'hC8;
	13'h865: q=8'hDE;
	13'h866: q=8'hF4;
	13'h867: q=8'hDF;
	13'h868: q=8'hAF;
	13'h869: q=8'hDE;
	13'h86A: q=8'hA5;
	13'h86B: q=8'hDF;
	13'h86C: q=8'hF4;
	13'h86D: q=8'hBD;
	13'h86E: q=8'h0;
	13'h86F: q=8'hF3;
	13'h870: q=8'h27;
	13'h871: q=8'h25;
	13'h872: q=8'hBD;
	13'h873: q=8'hEA;
	13'h874: q=8'h2F;
	13'h875: q=8'h20;
	13'h876: q=8'h9F;
	13'h877: q=8'hDF;
	13'h878: q=8'hF4;
	13'h879: q=8'hBD;
	13'h87A: q=8'hE6;
	13'h87B: q=8'h56;
	13'h87C: q=8'h8;
	13'h87D: q=8'h4D;
	13'h87E: q=8'h26;
	13'h87F: q=8'hF;
	13'h880: q=8'hC6;
	13'h881: q=8'h6;
	13'h882: q=8'hA6;
	13'h883: q=8'h0;
	13'h884: q=8'hAA;
	13'h885: q=8'h1;
	13'h886: q=8'h27;
	13'h887: q=8'h46;
	13'h888: q=8'hEC;
	13'h889: q=8'h2;
	13'h88A: q=8'hDD;
	13'h88B: q=8'hAB;
	13'h88C: q=8'hC6;
	13'h88D: q=8'h4;
	13'h88E: q=8'h3A;
	13'h88F: q=8'hA6;
	13'h890: q=8'h0;
	13'h891: q=8'h81;
	13'h892: q=8'h85;
	13'h893: q=8'h26;
	13'h894: q=8'hE2;
	13'h895: q=8'h20;
	13'h896: q=8'h97;
	13'h897: q=8'hDE;
	13'h898: q=8'hAF;
	13'h899: q=8'hD6;
	13'h89A: q=8'h87;
	13'h89B: q=8'h27;
	13'h89C: q=8'h3;
	13'h89D: q=8'h7E;
	13'h89E: q=8'hE5;
	13'h89F: q=8'h63;
	13'h8A0: q=8'hA6;
	13'h8A1: q=8'h0;
	13'h8A2: q=8'h27;
	13'h8A3: q=8'h6;
	13'h8A4: q=8'hCE;
	13'h8A5: q=8'hE8;
	13'h8A6: q=8'hAA;
	13'h8A7: q=8'h7E;
	13'h8A8: q=8'hE7;
	13'h8A9: q=8'hA8;
	13'h8AA: q=8'h39;
	13'h8AB: q=8'h3F;
	13'h8AC: q=8'h45;
	13'h8AD: q=8'h58;
	13'h8AE: q=8'h54;
	13'h8AF: q=8'h52;
	13'h8B0: q=8'h41;
	13'h8B1: q=8'h20;
	13'h8B2: q=8'h49;
	13'h8B3: q=8'h47;
	13'h8B4: q=8'h4E;
	13'h8B5: q=8'h4F;
	13'h8B6: q=8'h52;
	13'h8B7: q=8'h45;
	13'h8B8: q=8'h44;
	13'h8B9: q=8'hD;
	13'h8BA: q=8'h0;
	13'h8BB: q=8'h26;
	13'h8BC: q=8'h5;
	13'h8BD: q=8'hCE;
	13'h8BE: q=8'h0;
	13'h8BF: q=8'h0;
	13'h8C0: q=8'h20;
	13'h8C1: q=8'h3;
	13'h8C2: q=8'hBD;
	13'h8C3: q=8'hEB;
	13'h8C4: q=8'h1B;
	13'h8C5: q=8'hDF;
	13'h8C6: q=8'hB5;
	13'h8C7: q=8'hBD;
	13'h8C8: q=8'hE1;
	13'h8C9: q=8'hD8;
	13'h8CA: q=8'h27;
	13'h8CB: q=8'h4;
	13'h8CC: q=8'hC6;
	13'h8CD: q=8'h0;
	13'h8CE: q=8'h20;
	13'h8CF: q=8'h47;
	13'h8D0: q=8'h35;
	13'h8D1: q=8'h8;
	13'h8D2: q=8'h8;
	13'h8D3: q=8'h8;
	13'h8D4: q=8'hBD;
	13'h8D5: q=8'hF2;
	13'h8D6: q=8'h51;
	13'h8D7: q=8'h30;
	13'h8D8: q=8'hA6;
	13'h8D9: q=8'h8;
	13'h8DA: q=8'h97;
	13'h8DB: q=8'hCE;
	13'h8DC: q=8'hDE;
	13'h8DD: q=8'hB5;
	13'h8DE: q=8'hBD;
	13'h8DF: q=8'hEF;
	13'h8E0: q=8'h7D;
	13'h8E1: q=8'hBD;
	13'h8E2: q=8'hF2;
	13'h8E3: q=8'h70;
	13'h8E4: q=8'h30;
	13'h8E5: q=8'hC6;
	13'h8E6: q=8'h9;
	13'h8E7: q=8'h3A;
	13'h8E8: q=8'hBD;
	13'h8E9: q=8'hF2;
	13'h8EA: q=8'hD9;
	13'h8EB: q=8'h30;
	13'h8EC: q=8'hE0;
	13'h8ED: q=8'h8;
	13'h8EE: q=8'h27;
	13'h8EF: q=8'hC;
	13'h8F0: q=8'hEE;
	13'h8F1: q=8'hE;
	13'h8F2: q=8'hDF;
	13'h8F3: q=8'hE2;
	13'h8F4: q=8'h30;
	13'h8F5: q=8'hEE;
	13'h8F6: q=8'h10;
	13'h8F7: q=8'hDF;
	13'h8F8: q=8'hF4;
	13'h8F9: q=8'h7E;
	13'h8FA: q=8'hE5;
	13'h8FB: q=8'h19;
	13'h8FC: q=8'hC6;
	13'h8FD: q=8'h12;
	13'h8FE: q=8'h3A;
	13'h8FF: q=8'h35;
	13'h900: q=8'hBD;
	13'h901: q=8'h0;
	13'h902: q=8'hF3;
	13'h903: q=8'h81;
	13'h904: q=8'h2C;
	13'h905: q=8'h26;
	13'h906: q=8'hF2;
	13'h907: q=8'hBD;
	13'h908: q=8'h0;
	13'h909: q=8'hEB;
	13'h90A: q=8'h8D;
	13'h90B: q=8'hB6;
	13'h90C: q=8'h8D;
	13'h90D: q=8'hC;
	13'h90E: q=8'h6D;
	13'h90F: q=8'hD;
	13'h910: q=8'h76;
	13'h911: q=8'h0;
	13'h912: q=8'h84;
	13'h913: q=8'h28;
	13'h914: q=8'h95;
	13'h915: q=8'hC6;
	13'h916: q=8'h18;
	13'h917: q=8'h7E;
	13'h918: q=8'hE2;
	13'h919: q=8'h38;
	13'h91A: q=8'hDE;
	13'h91B: q=8'hF4;
	13'h91C: q=8'h9;
	13'h91D: q=8'hDF;
	13'h91E: q=8'hF4;
	13'h91F: q=8'h4F;
	13'h920: q=8'hC6;
	13'h921: q=8'h37;
	13'h922: q=8'h36;
	13'h923: q=8'hC6;
	13'h924: q=8'h1;
	13'h925: q=8'hBD;
	13'h926: q=8'hE2;
	13'h927: q=8'h1A;
	13'h928: q=8'hBD;
	13'h929: q=8'hE9;
	13'h92A: q=8'hE5;
	13'h92B: q=8'h7F;
	13'h92C: q=8'h0;
	13'h92D: q=8'hB9;
	13'h92E: q=8'hBD;
	13'h92F: q=8'h0;
	13'h930: q=8'hF3;
	13'h931: q=8'h80;
	13'h932: q=8'hAE;
	13'h933: q=8'h25;
	13'h934: q=8'h14;
	13'h935: q=8'h81;
	13'h936: q=8'h3;
	13'h937: q=8'h24;
	13'h938: q=8'h10;
	13'h939: q=8'h81;
	13'h93A: q=8'h1;
	13'h93B: q=8'h49;
	13'h93C: q=8'h98;
	13'h93D: q=8'hB9;
	13'h93E: q=8'h91;
	13'h93F: q=8'hB9;
	13'h940: q=8'h25;
	13'h941: q=8'h59;
	13'h942: q=8'h97;
	13'h943: q=8'hB9;
	13'h944: q=8'hBD;
	13'h945: q=8'h0;
	13'h946: q=8'hEB;
	13'h947: q=8'h20;
	13'h948: q=8'hE8;
	13'h949: q=8'hD6;
	13'h94A: q=8'hB9;
	13'h94B: q=8'h26;
	13'h94C: q=8'h2B;
	13'h94D: q=8'h24;
	13'h94E: q=8'h66;
	13'h94F: q=8'h8B;
	13'h950: q=8'h7;
	13'h951: q=8'h24;
	13'h952: q=8'h62;
	13'h953: q=8'h99;
	13'h954: q=8'h84;
	13'h955: q=8'h26;
	13'h956: q=8'h3;
	13'h957: q=8'h7E;
	13'h958: q=8'hEE;
	13'h959: q=8'h6;
	13'h95A: q=8'h89;
	13'h95B: q=8'hFF;
	13'h95C: q=8'h16;
	13'h95D: q=8'h48;
	13'h95E: q=8'h1B;
	13'h95F: q=8'h16;
	13'h960: q=8'hCE;
	13'h961: q=8'hE0;
	13'h962: q=8'h30;
	13'h963: q=8'h3A;
	13'h964: q=8'h32;
	13'h965: q=8'hA1;
	13'h966: q=8'h0;
	13'h967: q=8'h24;
	13'h968: q=8'h53;
	13'h969: q=8'h8D;
	13'h96A: q=8'hA3;
	13'h96B: q=8'h36;
	13'h96C: q=8'h8D;
	13'h96D: q=8'h23;
	13'h96E: q=8'hDE;
	13'h96F: q=8'hB7;
	13'h970: q=8'h32;
	13'h971: q=8'h26;
	13'h972: q=8'h18;
	13'h973: q=8'h4D;
	13'h974: q=8'h27;
	13'h975: q=8'h6C;
	13'h976: q=8'h20;
	13'h977: q=8'h4D;
	13'h978: q=8'h78;
	13'h979: q=8'h0;
	13'h97A: q=8'h84;
	13'h97B: q=8'h59;
	13'h97C: q=8'hDE;
	13'h97D: q=8'hF4;
	13'h97E: q=8'h9;
	13'h97F: q=8'hDF;
	13'h980: q=8'hF4;
	13'h981: q=8'hCE;
	13'h982: q=8'hE9;
	13'h983: q=8'h88;
	13'h984: q=8'hD7;
	13'h985: q=8'hB9;
	13'h986: q=8'h20;
	13'h987: q=8'hDC;
	13'h988: q=8'h64;
	13'h989: q=8'hEA;
	13'h98A: q=8'hAE;
	13'h98B: q=8'hA1;
	13'h98C: q=8'h0;
	13'h98D: q=8'h24;
	13'h98E: q=8'h36;
	13'h98F: q=8'h20;
	13'h990: q=8'hDA;
	13'h991: q=8'hEC;
	13'h992: q=8'h1;
	13'h993: q=8'h37;
	13'h994: q=8'h36;
	13'h995: q=8'h8D;
	13'h996: q=8'h7;
	13'h997: q=8'hD6;
	13'h998: q=8'hB9;
	13'h999: q=8'h20;
	13'h99A: q=8'h86;
	13'h99B: q=8'h7E;
	13'h99C: q=8'hEA;
	13'h99D: q=8'h3C;
	13'h99E: q=8'hD6;
	13'h99F: q=8'hCE;
	13'h9A0: q=8'hA6;
	13'h9A1: q=8'h0;
	13'h9A2: q=8'h38;
	13'h9A3: q=8'h37;
	13'h9A4: q=8'hD6;
	13'h9A5: q=8'hCD;
	13'h9A6: q=8'h37;
	13'h9A7: q=8'hD6;
	13'h9A8: q=8'hCC;
	13'h9A9: q=8'h37;
	13'h9AA: q=8'hD6;
	13'h9AB: q=8'hCB;
	13'h9AC: q=8'h37;
	13'h9AD: q=8'hD6;
	13'h9AE: q=8'hCA;
	13'h9AF: q=8'h37;
	13'h9B0: q=8'hD6;
	13'h9B1: q=8'hC9;
	13'h9B2: q=8'h37;
	13'h9B3: q=8'h6E;
	13'h9B4: q=8'h0;
	13'h9B5: q=8'hCE;
	13'h9B6: q=8'h0;
	13'h9B7: q=8'h0;
	13'h9B8: q=8'h32;
	13'h9B9: q=8'h4D;
	13'h9BA: q=8'h27;
	13'h9BB: q=8'h26;
	13'h9BC: q=8'h81;
	13'h9BD: q=8'h64;
	13'h9BE: q=8'h27;
	13'h9BF: q=8'h3;
	13'h9C0: q=8'hBD;
	13'h9C1: q=8'hE9;
	13'h9C2: q=8'hE;
	13'h9C3: q=8'hDF;
	13'h9C4: q=8'hB7;
	13'h9C5: q=8'h33;
	13'h9C6: q=8'h81;
	13'h9C7: q=8'h5A;
	13'h9C8: q=8'h27;
	13'h9C9: q=8'h1A;
	13'h9CA: q=8'h81;
	13'h9CB: q=8'h7D;
	13'h9CC: q=8'h27;
	13'h9CD: q=8'h16;
	13'h9CE: q=8'h54;
	13'h9CF: q=8'hD7;
	13'h9D0: q=8'h88;
	13'h9D1: q=8'h32;
	13'h9D2: q=8'h33;
	13'h9D3: q=8'hDD;
	13'h9D4: q=8'hD6;
	13'h9D5: q=8'h38;
	13'h9D6: q=8'hDF;
	13'h9D7: q=8'hD8;
	13'h9D8: q=8'h33;
	13'h9D9: q=8'hD7;
	13'h9DA: q=8'hDA;
	13'h9DB: q=8'h33;
	13'h9DC: q=8'hD7;
	13'h9DD: q=8'hDB;
	13'h9DE: q=8'hD8;
	13'h9DF: q=8'hCE;
	13'h9E0: q=8'hD7;
	13'h9E1: q=8'hDC;
	13'h9E2: q=8'hD6;
	13'h9E3: q=8'hC9;
	13'h9E4: q=8'h39;
	13'h9E5: q=8'hBD;
	13'h9E6: q=8'h42;
	13'h9E7: q=8'h94;
	13'h9E8: q=8'h7F;
	13'h9E9: q=8'h0;
	13'h9EA: q=8'h84;
	13'h9EB: q=8'h8D;
	13'h9EC: q=8'h4C;
	13'h9ED: q=8'h24;
	13'h9EE: q=8'h3;
	13'h9EF: q=8'h7E;
	13'h9F0: q=8'hF3;
	13'h9F1: q=8'h59;
	13'h9F2: q=8'hBD;
	13'h9F3: q=8'hEB;
	13'h9F4: q=8'h76;
	13'h9F5: q=8'h24;
	13'h9F6: q=8'h52;
	13'h9F7: q=8'h81;
	13'h9F8: q=8'h2E;
	13'h9F9: q=8'h27;
	13'h9FA: q=8'hF4;
	13'h9FB: q=8'h81;
	13'h9FC: q=8'hA8;
	13'h9FD: q=8'h27;
	13'h9FE: q=8'h42;
	13'h9FF: q=8'h81;
	13'hA00: q=8'hA7;
	13'hA01: q=8'h27;
	13'hA02: q=8'hE2;
	13'hA03: q=8'h81;
	13'hA04: q=8'h22;
	13'hA05: q=8'h26;
	13'hA06: q=8'h8;
	13'hA07: q=8'hDE;
	13'hA08: q=8'hF4;
	13'hA09: q=8'hBD;
	13'hA0A: q=8'hED;
	13'hA0B: q=8'h6;
	13'hA0C: q=8'h7E;
	13'hA0D: q=8'hEF;
	13'hA0E: q=8'h3E;
	13'hA0F: q=8'h81;
	13'hA10: q=8'hA4;
	13'hA11: q=8'h26;
	13'hA12: q=8'hD;
	13'hA13: q=8'h86;
	13'hA14: q=8'h5A;
	13'hA15: q=8'hBD;
	13'hA16: q=8'hE9;
	13'hA17: q=8'h21;
	13'hA18: q=8'hBD;
	13'hA19: q=8'hEB;
	13'hA1A: q=8'hC7;
	13'hA1B: q=8'h43;
	13'hA1C: q=8'h53;
	13'hA1D: q=8'h7E;
	13'hA1E: q=8'hEC;
	13'hA1F: q=8'hE3;
	13'hA20: q=8'h80;
	13'hA21: q=8'hB1;
	13'hA22: q=8'h24;
	13'hA23: q=8'h31;
	13'hA24: q=8'h8D;
	13'hA25: q=8'h6;
	13'hA26: q=8'hBD;
	13'hA27: q=8'hE9;
	13'hA28: q=8'h1A;
	13'hA29: q=8'hC6;
	13'hA2A: q=8'h29;
	13'hA2B: q=8'h8C;
	13'hA2C: q=8'hC6;
	13'hA2D: q=8'h28;
	13'hA2E: q=8'h8C;
	13'hA2F: q=8'hC6;
	13'hA30: q=8'h2C;
	13'hA31: q=8'h3C;
	13'hA32: q=8'hDE;
	13'hA33: q=8'hF4;
	13'hA34: q=8'hE1;
	13'hA35: q=8'h0;
	13'hA36: q=8'h38;
	13'hA37: q=8'h26;
	13'hA38: q=8'h3;
	13'hA39: q=8'h7E;
	13'hA3A: q=8'h0;
	13'hA3B: q=8'hEB;
	13'hA3C: q=8'hC6;
	13'hA3D: q=8'h2;
	13'hA3E: q=8'h7E;
	13'hA3F: q=8'hE2;
	13'hA40: q=8'h38;
	13'hA41: q=8'h86;
	13'hA42: q=8'h7D;
	13'hA43: q=8'hBD;
	13'hA44: q=8'hE9;
	13'hA45: q=8'h21;
	13'hA46: q=8'h7E;
	13'hA47: q=8'hF5;
	13'hA48: q=8'h93;
	13'hA49: q=8'hBD;
	13'hA4A: q=8'hEB;
	13'hA4B: q=8'h1B;
	13'hA4C: q=8'hDF;
	13'hA4D: q=8'hCC;
	13'hA4E: q=8'h96;
	13'hA4F: q=8'h84;
	13'hA50: q=8'h26;
	13'hA51: q=8'h92;
	13'hA52: q=8'h7E;
	13'hA53: q=8'hF2;
	13'hA54: q=8'h51;
	13'hA55: q=8'h16;
	13'hA56: q=8'h58;
	13'hA57: q=8'h8D;
	13'hA58: q=8'hE0;
	13'hA59: q=8'h37;
	13'hA5A: q=8'hC1;
	13'hA5B: q=8'h22;
	13'hA5C: q=8'h25;
	13'hA5D: q=8'h21;
	13'hA5E: q=8'hC1;
	13'hA5F: q=8'h2C;
	13'hA60: q=8'h24;
	13'hA61: q=8'h1F;
	13'hA62: q=8'h8D;
	13'hA63: q=8'hC8;
	13'hA64: q=8'h33;
	13'hA65: q=8'hC1;
	13'hA66: q=8'h28;
	13'hA67: q=8'h24;
	13'hA68: q=8'h19;
	13'hA69: q=8'h37;
	13'hA6A: q=8'hBD;
	13'hA6B: q=8'hE9;
	13'hA6C: q=8'h1A;
	13'hA6D: q=8'h8D;
	13'hA6E: q=8'hC0;
	13'hA6F: q=8'hBD;
	13'hA70: q=8'hE9;
	13'hA71: q=8'hF;
	13'hA72: q=8'h32;
	13'hA73: q=8'hDE;
	13'hA74: q=8'hCC;
	13'hA75: q=8'h3C;
	13'hA76: q=8'h36;
	13'hA77: q=8'hBD;
	13'hA78: q=8'hEF;
	13'hA79: q=8'hD;
	13'hA7A: q=8'h32;
	13'hA7B: q=8'h37;
	13'hA7C: q=8'h16;
	13'hA7D: q=8'h20;
	13'hA7E: q=8'h3;
	13'hA7F: q=8'h8D;
	13'hA80: q=8'hA3;
	13'hA81: q=8'h33;
	13'hA82: q=8'hCE;
	13'hA83: q=8'hE0;
	13'hA84: q=8'h0;
	13'hA85: q=8'h3A;
	13'hA86: q=8'hEE;
	13'hA87: q=8'h0;
	13'hA88: q=8'hAD;
	13'hA89: q=8'h0;
	13'hA8A: q=8'h7E;
	13'hA8B: q=8'hE9;
	13'hA8C: q=8'hE;
	13'hA8D: q=8'h86;
	13'hA8E: q=8'h4F;
	13'hA8F: q=8'h97;
	13'hA90: q=8'h82;
	13'hA91: q=8'hBD;
	13'hA92: q=8'hEB;
	13'hA93: q=8'hC7;
	13'hA94: q=8'hDD;
	13'hA95: q=8'h80;
	13'hA96: q=8'hBD;
	13'hA97: q=8'hF2;
	13'hA98: q=8'h8B;
	13'hA99: q=8'hBD;
	13'hA9A: q=8'hEB;
	13'hA9B: q=8'hC7;
	13'hA9C: q=8'h7D;
	13'hA9D: q=8'h0;
	13'hA9E: q=8'h82;
	13'hA9F: q=8'h26;
	13'hAA0: q=8'h6;
	13'hAA1: q=8'h94;
	13'hAA2: q=8'h80;
	13'hAA3: q=8'hD4;
	13'hAA4: q=8'h81;
	13'hAA5: q=8'h20;
	13'hAA6: q=8'h4;
	13'hAA7: q=8'h9A;
	13'hAA8: q=8'h80;
	13'hAA9: q=8'hDA;
	13'hAAA: q=8'h81;
	13'hAAB: q=8'h7E;
	13'hAAC: q=8'hEC;
	13'hAAD: q=8'hE3;
	13'hAAE: q=8'hBD;
	13'hAAF: q=8'hE9;
	13'hAB0: q=8'h10;
	13'hAB1: q=8'h26;
	13'hAB2: q=8'h10;
	13'hAB3: q=8'h96;
	13'hAB4: q=8'hDB;
	13'hAB5: q=8'h8A;
	13'hAB6: q=8'h7F;
	13'hAB7: q=8'h94;
	13'hAB8: q=8'hD7;
	13'hAB9: q=8'h97;
	13'hABA: q=8'hD7;
	13'hABB: q=8'hCE;
	13'hABC: q=8'h0;
	13'hABD: q=8'hD6;
	13'hABE: q=8'hBD;
	13'hABF: q=8'hF2;
	13'hAC0: q=8'hD9;
	13'hAC1: q=8'h20;
	13'hAC2: q=8'h40;
	13'hAC3: q=8'h7F;
	13'hAC4: q=8'h0;
	13'hAC5: q=8'h84;
	13'hAC6: q=8'h7A;
	13'hAC7: q=8'h0;
	13'hAC8: q=8'hB9;
	13'hAC9: q=8'hBD;
	13'hACA: q=8'hEE;
	13'hACB: q=8'h56;
	13'hACC: q=8'hD7;
	13'hACD: q=8'hD0;
	13'hACE: q=8'hDF;
	13'hACF: q=8'hD2;
	13'hAD0: q=8'hDE;
	13'hAD1: q=8'hD9;
	13'hAD2: q=8'hBD;
	13'hAD3: q=8'hEE;
	13'hAD4: q=8'h58;
	13'hAD5: q=8'h96;
	13'hAD6: q=8'hD0;
	13'hAD7: q=8'h10;
	13'hAD8: q=8'h27;
	13'hAD9: q=8'h7;
	13'hADA: q=8'h86;
	13'hADB: q=8'h1;
	13'hADC: q=8'h24;
	13'hADD: q=8'h3;
	13'hADE: q=8'hD6;
	13'hADF: q=8'hD0;
	13'hAE0: q=8'h40;
	13'hAE1: q=8'h97;
	13'hAE2: q=8'hCE;
	13'hAE3: q=8'h7;
	13'hAE4: q=8'h36;
	13'hAE5: q=8'h9F;
	13'hAE6: q=8'h91;
	13'hAE7: q=8'hF;
	13'hAE8: q=8'h35;
	13'hAE9: q=8'hDE;
	13'hAEA: q=8'hD2;
	13'hAEB: q=8'h5C;
	13'hAEC: q=8'h9;
	13'hAED: q=8'h5A;
	13'hAEE: q=8'h26;
	13'hAEF: q=8'h4;
	13'hAF0: q=8'hD6;
	13'hAF1: q=8'hCE;
	13'hAF2: q=8'h20;
	13'hAF3: q=8'hB;
	13'hAF4: q=8'h32;
	13'hAF5: q=8'h8;
	13'hAF6: q=8'hA1;
	13'hAF7: q=8'h0;
	13'hAF8: q=8'h27;
	13'hAF9: q=8'hF3;
	13'hAFA: q=8'hC6;
	13'hAFB: q=8'hFF;
	13'hAFC: q=8'h24;
	13'hAFD: q=8'h1;
	13'hAFE: q=8'h50;
	13'hAFF: q=8'h9E;
	13'hB00: q=8'h91;
	13'hB01: q=8'h32;
	13'hB02: q=8'h6;
	13'hB03: q=8'hCB;
	13'hB04: q=8'h1;
	13'hB05: q=8'h59;
	13'hB06: q=8'hD4;
	13'hB07: q=8'h88;
	13'hB08: q=8'h27;
	13'hB09: q=8'h2;
	13'hB0A: q=8'hC6;
	13'hB0B: q=8'hFF;
	13'hB0C: q=8'h7E;
	13'hB0D: q=8'hF2;
	13'hB0E: q=8'hBC;
	13'hB0F: q=8'hBD;
	13'hB10: q=8'hEA;
	13'hB11: q=8'h2F;
	13'hB12: q=8'h16;
	13'hB13: q=8'h8D;
	13'hB14: q=8'hA;
	13'hB15: q=8'hBD;
	13'hB16: q=8'h0;
	13'hB17: q=8'hF3;
	13'hB18: q=8'h26;
	13'hB19: q=8'hF5;
	13'hB1A: q=8'h39;
	13'hB1B: q=8'h5F;
	13'hB1C: q=8'hBD;
	13'hB1D: q=8'h0;
	13'hB1E: q=8'hF3;
	13'hB1F: q=8'hD7;
	13'hB20: q=8'h83;
	13'hB21: q=8'h97;
	13'hB22: q=8'hB1;
	13'hB23: q=8'hBD;
	13'hB24: q=8'h0;
	13'hB25: q=8'hF3;
	13'hB26: q=8'h8D;
	13'hB27: q=8'h4E;
	13'hB28: q=8'h24;
	13'hB29: q=8'h3;
	13'hB2A: q=8'h7E;
	13'hB2B: q=8'hEA;
	13'hB2C: q=8'h3C;
	13'hB2D: q=8'h5F;
	13'hB2E: q=8'hD7;
	13'hB2F: q=8'h84;
	13'hB30: q=8'hBD;
	13'hB31: q=8'h0;
	13'hB32: q=8'hEB;
	13'hB33: q=8'h25;
	13'hB34: q=8'h4;
	13'hB35: q=8'h8D;
	13'hB36: q=8'h3F;
	13'hB37: q=8'h25;
	13'hB38: q=8'hA;
	13'hB39: q=8'h16;
	13'hB3A: q=8'hBD;
	13'hB3B: q=8'h0;
	13'hB3C: q=8'hEB;
	13'hB3D: q=8'h25;
	13'hB3E: q=8'hFB;
	13'hB3F: q=8'h8D;
	13'hB40: q=8'h35;
	13'hB41: q=8'h24;
	13'hB42: q=8'hF7;
	13'hB43: q=8'h81;
	13'hB44: q=8'h24;
	13'hB45: q=8'h26;
	13'hB46: q=8'h8;
	13'hB47: q=8'h73;
	13'hB48: q=8'h0;
	13'hB49: q=8'h84;
	13'hB4A: q=8'hCB;
	13'hB4B: q=8'h80;
	13'hB4C: q=8'hBD;
	13'hB4D: q=8'h0;
	13'hB4E: q=8'hEB;
	13'hB4F: q=8'hD7;
	13'hB50: q=8'hB2;
	13'hB51: q=8'hD6;
	13'hB52: q=8'h86;
	13'hB53: q=8'h5A;
	13'hB54: q=8'h26;
	13'hB55: q=8'h3;
	13'hB56: q=8'h7E;
	13'hB57: q=8'hEC;
	13'hB58: q=8'h7;
	13'hB59: q=8'h9B;
	13'hB5A: q=8'h86;
	13'hB5B: q=8'h80;
	13'hB5C: q=8'h28;
	13'hB5D: q=8'h26;
	13'hB5E: q=8'h3;
	13'hB5F: q=8'h7E;
	13'hB60: q=8'hEB;
	13'hB61: q=8'hDE;
	13'hB62: q=8'h7F;
	13'hB63: q=8'h0;
	13'hB64: q=8'h86;
	13'hB65: q=8'hDE;
	13'hB66: q=8'h95;
	13'hB67: q=8'h9C;
	13'hB68: q=8'h97;
	13'hB69: q=8'h27;
	13'hB6A: q=8'h14;
	13'hB6B: q=8'hDC;
	13'hB6C: q=8'hB1;
	13'hB6D: q=8'hA3;
	13'hB6E: q=8'h0;
	13'hB6F: q=8'h27;
	13'hB70: q=8'h3F;
	13'hB71: q=8'hC6;
	13'hB72: q=8'h7;
	13'hB73: q=8'h3A;
	13'hB74: q=8'h20;
	13'hB75: q=8'hF1;
	13'hB76: q=8'h81;
	13'hB77: q=8'h41;
	13'hB78: q=8'h25;
	13'hB79: q=8'h4;
	13'hB7A: q=8'h80;
	13'hB7B: q=8'h5B;
	13'hB7C: q=8'h80;
	13'hB7D: q=8'hA5;
	13'hB7E: q=8'h39;
	13'hB7F: q=8'h38;
	13'hB80: q=8'h3C;
	13'hB81: q=8'h8C;
	13'hB82: q=8'hEA;
	13'hB83: q=8'h4C;
	13'hB84: q=8'h26;
	13'hB85: q=8'h4;
	13'hB86: q=8'hCE;
	13'hB87: q=8'hEB;
	13'hB88: q=8'hB7;
	13'hB89: q=8'h39;
	13'hB8A: q=8'hDC;
	13'hB8B: q=8'h99;
	13'hB8C: q=8'hDD;
	13'hB8D: q=8'hBD;
	13'hB8E: q=8'hC3;
	13'hB8F: q=8'h0;
	13'hB90: q=8'h7;
	13'hB91: q=8'hDD;
	13'hB92: q=8'hBB;
	13'hB93: q=8'hDE;
	13'hB94: q=8'h97;
	13'hB95: q=8'hDF;
	13'hB96: q=8'hC1;
	13'hB97: q=8'hBD;
	13'hB98: q=8'hE1;
	13'hB99: q=8'hFE;
	13'hB9A: q=8'hDE;
	13'hB9B: q=8'hBB;
	13'hB9C: q=8'hDF;
	13'hB9D: q=8'h99;
	13'hB9E: q=8'hDE;
	13'hB9F: q=8'hBF;
	13'hBA0: q=8'hDF;
	13'hBA1: q=8'h97;
	13'hBA2: q=8'hDE;
	13'hBA3: q=8'hC1;
	13'hBA4: q=8'hDC;
	13'hBA5: q=8'hB1;
	13'hBA6: q=8'hED;
	13'hBA7: q=8'h0;
	13'hBA8: q=8'h4F;
	13'hBA9: q=8'h5F;
	13'hBAA: q=8'hED;
	13'hBAB: q=8'h2;
	13'hBAC: q=8'hED;
	13'hBAD: q=8'h4;
	13'hBAE: q=8'hA7;
	13'hBAF: q=8'h6;
	13'hBB0: q=8'h8;
	13'hBB1: q=8'h8;
	13'hBB2: q=8'hDF;
	13'hBB3: q=8'hB3;
	13'hBB4: q=8'h39;
	13'hBB5: q=8'h90;
	13'hBB6: q=8'h80;
	13'hBB7: q=8'h0;
	13'hBB8: q=8'h0;
	13'hBB9: q=8'h0;
	13'hBBA: q=8'hBD;
	13'hBBB: q=8'h0;
	13'hBBC: q=8'hEB;
	13'hBBD: q=8'hBD;
	13'hBBE: q=8'hE9;
	13'hBBF: q=8'hC;
	13'hBC0: q=8'hBD;
	13'hBC1: q=8'hE9;
	13'hBC2: q=8'hE;
	13'hBC3: q=8'h96;
	13'hBC4: q=8'hCE;
	13'hBC5: q=8'h2B;
	13'hBC6: q=8'h67;
	13'hBC7: q=8'hBD;
	13'hBC8: q=8'hE9;
	13'hBC9: q=8'hE;
	13'hBCA: q=8'h96;
	13'hBCB: q=8'hC9;
	13'hBCC: q=8'h81;
	13'hBCD: q=8'h90;
	13'hBCE: q=8'h25;
	13'hBCF: q=8'h8;
	13'hBD0: q=8'hCE;
	13'hBD1: q=8'hEB;
	13'hBD2: q=8'hB5;
	13'hBD3: q=8'hBD;
	13'hBD4: q=8'hF2;
	13'hBD5: q=8'hD9;
	13'hBD6: q=8'h26;
	13'hBD7: q=8'h56;
	13'hBD8: q=8'hBD;
	13'hBD9: q=8'hF3;
	13'hBDA: q=8'hB;
	13'hBDB: q=8'hDC;
	13'hBDC: q=8'hCC;
	13'hBDD: q=8'h39;
	13'hBDE: q=8'hDE;
	13'hBDF: q=8'h83;
	13'hBE0: q=8'h3C;
	13'hBE1: q=8'h5F;
	13'hBE2: q=8'h37;
	13'hBE3: q=8'hDE;
	13'hBE4: q=8'hB1;
	13'hBE5: q=8'h3C;
	13'hBE6: q=8'h8D;
	13'hBE7: q=8'hD2;
	13'hBE8: q=8'h38;
	13'hBE9: q=8'hDF;
	13'hBEA: q=8'hB1;
	13'hBEB: q=8'h33;
	13'hBEC: q=8'h5C;
	13'hBED: q=8'hD7;
	13'hBEE: q=8'h82;
	13'hBEF: q=8'h32;
	13'hBF0: q=8'h33;
	13'hBF1: q=8'hDE;
	13'hBF2: q=8'hCC;
	13'hBF3: q=8'h3C;
	13'hBF4: q=8'h37;
	13'hBF5: q=8'h36;
	13'hBF6: q=8'hD6;
	13'hBF7: q=8'h82;
	13'hBF8: q=8'hBD;
	13'hBF9: q=8'h0;
	13'hBFA: q=8'hF3;
	13'hBFB: q=8'h81;
	13'hBFC: q=8'h2C;
	13'hBFD: q=8'h27;
	13'hBFE: q=8'hE3;
	13'hBFF: q=8'hBD;
	13'hC00: q=8'hEA;
	13'hC01: q=8'h29;
	13'hC02: q=8'h38;
	13'hC03: q=8'hDF;
	13'hC04: q=8'h83;
	13'hC05: q=8'hC6;
	13'hC06: q=8'hFF;
	13'hC07: q=8'h37;
	13'hC08: q=8'hDE;
	13'hC09: q=8'h97;
	13'hC0A: q=8'h9C;
	13'hC0B: q=8'h99;
	13'hC0C: q=8'h27;
	13'hC0D: q=8'h25;
	13'hC0E: q=8'hDC;
	13'hC0F: q=8'hB1;
	13'hC10: q=8'hA3;
	13'hC11: q=8'h0;
	13'hC12: q=8'h27;
	13'hC13: q=8'h7;
	13'hC14: q=8'hEC;
	13'hC15: q=8'h2;
	13'hC16: q=8'hBD;
	13'hC17: q=8'hE2;
	13'hC18: q=8'h2D;
	13'hC19: q=8'h20;
	13'hC1A: q=8'hEF;
	13'hC1B: q=8'hC6;
	13'hC1C: q=8'h12;
	13'hC1D: q=8'h32;
	13'hC1E: q=8'h4D;
	13'hC1F: q=8'h27;
	13'hC20: q=8'hBC;
	13'hC21: q=8'h96;
	13'hC22: q=8'h83;
	13'hC23: q=8'h26;
	13'hC24: q=8'hB;
	13'hC25: q=8'hD6;
	13'hC26: q=8'h82;
	13'hC27: q=8'hE1;
	13'hC28: q=8'h4;
	13'hC29: q=8'h27;
	13'hC2A: q=8'h5C;
	13'hC2B: q=8'hC6;
	13'hC2C: q=8'h10;
	13'hC2D: q=8'h8C;
	13'hC2E: q=8'hC6;
	13'hC2F: q=8'h8;
	13'hC30: q=8'h7E;
	13'hC31: q=8'hE2;
	13'hC32: q=8'h38;
	13'hC33: q=8'h32;
	13'hC34: q=8'h4D;
	13'hC35: q=8'h27;
	13'hC36: q=8'hF7;
	13'hC37: q=8'hCC;
	13'hC38: q=8'h0;
	13'hC39: q=8'h5;
	13'hC3A: q=8'hDD;
	13'hC3B: q=8'hDE;
	13'hC3C: q=8'hDC;
	13'hC3D: q=8'hB1;
	13'hC3E: q=8'hED;
	13'hC3F: q=8'h0;
	13'hC40: q=8'hD6;
	13'hC41: q=8'h82;
	13'hC42: q=8'hE7;
	13'hC43: q=8'h4;
	13'hC44: q=8'hBD;
	13'hC45: q=8'hE2;
	13'hC46: q=8'h1A;
	13'hC47: q=8'hDF;
	13'hC48: q=8'hBB;
	13'hC49: q=8'hC6;
	13'hC4A: q=8'hB;
	13'hC4B: q=8'h4F;
	13'hC4C: q=8'h7D;
	13'hC4D: q=8'h0;
	13'hC4E: q=8'h83;
	13'hC4F: q=8'h27;
	13'hC50: q=8'h5;
	13'hC51: q=8'h32;
	13'hC52: q=8'h33;
	13'hC53: q=8'hC3;
	13'hC54: q=8'h0;
	13'hC55: q=8'h1;
	13'hC56: q=8'hED;
	13'hC57: q=8'h5;
	13'hC58: q=8'h8D;
	13'hC59: q=8'h5F;
	13'hC5A: q=8'hDD;
	13'hC5B: q=8'hDE;
	13'hC5C: q=8'h8;
	13'hC5D: q=8'h8;
	13'hC5E: q=8'h7A;
	13'hC5F: q=8'h0;
	13'hC60: q=8'h82;
	13'hC61: q=8'h26;
	13'hC62: q=8'hE6;
	13'hC63: q=8'hBD;
	13'hC64: q=8'hE2;
	13'hC65: q=8'h2D;
	13'hC66: q=8'h24;
	13'hC67: q=8'h3;
	13'hC68: q=8'h7E;
	13'hC69: q=8'hE2;
	13'hC6A: q=8'h36;
	13'hC6B: q=8'hBD;
	13'hC6C: q=8'hE2;
	13'hC6D: q=8'h1E;
	13'hC6E: q=8'h83;
	13'hC6F: q=8'h0;
	13'hC70: q=8'h35;
	13'hC71: q=8'hDD;
	13'hC72: q=8'h99;
	13'hC73: q=8'h4F;
	13'hC74: q=8'h9;
	13'hC75: q=8'hA7;
	13'hC76: q=8'h5;
	13'hC77: q=8'h9C;
	13'hC78: q=8'h89;
	13'hC79: q=8'h26;
	13'hC7A: q=8'hF9;
	13'hC7B: q=8'hDE;
	13'hC7C: q=8'hBB;
	13'hC7D: q=8'h96;
	13'hC7E: q=8'h99;
	13'hC7F: q=8'h93;
	13'hC80: q=8'hBB;
	13'hC81: q=8'hED;
	13'hC82: q=8'h2;
	13'hC83: q=8'h96;
	13'hC84: q=8'h83;
	13'hC85: q=8'h26;
	13'hC86: q=8'h31;
	13'hC87: q=8'hE6;
	13'hC88: q=8'h4;
	13'hC89: q=8'hD7;
	13'hC8A: q=8'h82;
	13'hC8B: q=8'h4F;
	13'hC8C: q=8'h5F;
	13'hC8D: q=8'hDD;
	13'hC8E: q=8'hDE;
	13'hC8F: q=8'h32;
	13'hC90: q=8'h33;
	13'hC91: q=8'hDD;
	13'hC92: q=8'hCC;
	13'hC93: q=8'h37;
	13'hC94: q=8'h36;
	13'hC95: q=8'hA3;
	13'hC96: q=8'h5;
	13'hC97: q=8'h24;
	13'hC98: q=8'h3F;
	13'hC99: q=8'hDC;
	13'hC9A: q=8'hDE;
	13'hC9B: q=8'h32;
	13'hC9C: q=8'h33;
	13'hC9D: q=8'h27;
	13'hC9E: q=8'h4;
	13'hC9F: q=8'h8D;
	13'hCA0: q=8'h18;
	13'hCA1: q=8'hD3;
	13'hCA2: q=8'hCC;
	13'hCA3: q=8'h8;
	13'hCA4: q=8'h8;
	13'hCA5: q=8'h7A;
	13'hCA6: q=8'h0;
	13'hCA7: q=8'h82;
	13'hCA8: q=8'h26;
	13'hCA9: q=8'hE3;
	13'hCAA: q=8'hDD;
	13'hCAB: q=8'h89;
	13'hCAC: q=8'h5;
	13'hCAD: q=8'h5;
	13'hCAE: q=8'hD3;
	13'hCAF: q=8'h89;
	13'hCB0: q=8'hC3;
	13'hCB1: q=8'h0;
	13'hCB2: q=8'h5;
	13'hCB3: q=8'hBD;
	13'hCB4: q=8'hE2;
	13'hCB5: q=8'h2D;
	13'hCB6: q=8'hDF;
	13'hCB7: q=8'hB3;
	13'hCB8: q=8'h39;
	13'hCB9: q=8'h86;
	13'hCBA: q=8'h10;
	13'hCBB: q=8'h97;
	13'hCBC: q=8'hBF;
	13'hCBD: q=8'hEC;
	13'hCBE: q=8'h5;
	13'hCBF: q=8'hDD;
	13'hCC0: q=8'h91;
	13'hCC1: q=8'h4F;
	13'hCC2: q=8'h5F;
	13'hCC3: q=8'h5;
	13'hCC4: q=8'h25;
	13'hCC5: q=8'h12;
	13'hCC6: q=8'h78;
	13'hCC7: q=8'h0;
	13'hCC8: q=8'hDF;
	13'hCC9: q=8'h79;
	13'hCCA: q=8'h0;
	13'hCCB: q=8'hDE;
	13'hCCC: q=8'h24;
	13'hCCD: q=8'h4;
	13'hCCE: q=8'hD3;
	13'hCCF: q=8'h91;
	13'hCD0: q=8'h25;
	13'hCD1: q=8'h6;
	13'hCD2: q=8'h7A;
	13'hCD3: q=8'h0;
	13'hCD4: q=8'hBF;
	13'hCD5: q=8'h26;
	13'hCD6: q=8'hEC;
	13'hCD7: q=8'h39;
	13'hCD8: q=8'h7E;
	13'hCD9: q=8'hEC;
	13'hCDA: q=8'h2B;
	13'hCDB: q=8'h9F;
	13'hCDC: q=8'h91;
	13'hCDD: q=8'hDC;
	13'hCDE: q=8'h91;
	13'hCDF: q=8'h93;
	13'hCE0: q=8'h99;
	13'hCE1: q=8'h21;
	13'hCE2: q=8'h4F;
	13'hCE3: q=8'h7F;
	13'hCE4: q=8'h0;
	13'hCE5: q=8'h84;
	13'hCE6: q=8'hDD;
	13'hCE7: q=8'hCA;
	13'hCE8: q=8'hC6;
	13'hCE9: q=8'h90;
	13'hCEA: q=8'h7E;
	13'hCEB: q=8'hF2;
	13'hCEC: q=8'hC3;
	13'hCED: q=8'hBD;
	13'hCEE: q=8'hE9;
	13'hCEF: q=8'hE;
	13'hCF0: q=8'hCE;
	13'hCF1: q=8'h43;
	13'hCF2: q=8'h34;
	13'hCF3: q=8'hBD;
	13'hCF4: q=8'hF4;
	13'hCF5: q=8'h29;
	13'hCF6: q=8'h38;
	13'hCF7: q=8'hCE;
	13'hCF8: q=8'h43;
	13'hCF9: q=8'h33;
	13'hCFA: q=8'h20;
	13'hCFB: q=8'hA;
	13'hCFC: q=8'hDF;
	13'hCFD: q=8'hC7;
	13'hCFE: q=8'h8D;
	13'hCFF: q=8'h5F;
	13'hD00: q=8'hDF;
	13'hD01: q=8'hD2;
	13'hD02: q=8'hD7;
	13'hD03: q=8'hD0;
	13'hD04: q=8'h39;
	13'hD05: q=8'h9;
	13'hD06: q=8'h86;
	13'hD07: q=8'h22;
	13'hD08: q=8'h97;
	13'hD09: q=8'h80;
	13'hD0A: q=8'h97;
	13'hD0B: q=8'h81;
	13'hD0C: q=8'h8;
	13'hD0D: q=8'hDF;
	13'hD0E: q=8'hDC;
	13'hD0F: q=8'hDF;
	13'hD10: q=8'hD2;
	13'hD11: q=8'hC6;
	13'hD12: q=8'hFF;
	13'hD13: q=8'h5C;
	13'hD14: q=8'hA6;
	13'hD15: q=8'h0;
	13'hD16: q=8'h27;
	13'hD17: q=8'hE;
	13'hD18: q=8'h8;
	13'hD19: q=8'h91;
	13'hD1A: q=8'h80;
	13'hD1B: q=8'h27;
	13'hD1C: q=8'h4;
	13'hD1D: q=8'h91;
	13'hD1E: q=8'h81;
	13'hD1F: q=8'h26;
	13'hD20: q=8'hF2;
	13'hD21: q=8'h81;
	13'hD22: q=8'h22;
	13'hD23: q=8'h27;
	13'hD24: q=8'h1;
	13'hD25: q=8'h9;
	13'hD26: q=8'hDF;
	13'hD27: q=8'hDE;
	13'hD28: q=8'hD7;
	13'hD29: q=8'hD0;
	13'hD2A: q=8'h37;
	13'hD2B: q=8'hDC;
	13'hD2C: q=8'hDC;
	13'hD2D: q=8'h83;
	13'hD2E: q=8'h43;
	13'hD2F: q=8'h34;
	13'hD30: q=8'h33;
	13'hD31: q=8'h22;
	13'hD32: q=8'h7;
	13'hD33: q=8'h8D;
	13'hD34: q=8'hC7;
	13'hD35: q=8'hDE;
	13'hD36: q=8'hDC;
	13'hD37: q=8'hBD;
	13'hD38: q=8'hEE;
	13'hD39: q=8'h3A;
	13'hD3A: q=8'hFE;
	13'hD3B: q=8'h42;
	13'hD3C: q=8'h3D;
	13'hD3D: q=8'h8C;
	13'hD3E: q=8'h42;
	13'hD3F: q=8'h50;
	13'hD40: q=8'h26;
	13'hD41: q=8'h5;
	13'hD42: q=8'hC6;
	13'hD43: q=8'h1E;
	13'hD44: q=8'h7E;
	13'hD45: q=8'hE2;
	13'hD46: q=8'h38;
	13'hD47: q=8'h96;
	13'hD48: q=8'hD0;
	13'hD49: q=8'hA7;
	13'hD4A: q=8'h0;
	13'hD4B: q=8'hDC;
	13'hD4C: q=8'hD2;
	13'hD4D: q=8'hED;
	13'hD4E: q=8'h2;
	13'hD4F: q=8'h86;
	13'hD50: q=8'hFF;
	13'hD51: q=8'h97;
	13'hD52: q=8'h84;
	13'hD53: q=8'hFF;
	13'hD54: q=8'h42;
	13'hD55: q=8'h3F;
	13'hD56: q=8'hDF;
	13'hD57: q=8'hCC;
	13'hD58: q=8'hC6;
	13'hD59: q=8'h5;
	13'hD5A: q=8'h3A;
	13'hD5B: q=8'hFF;
	13'hD5C: q=8'h42;
	13'hD5D: q=8'h3D;
	13'hD5E: q=8'h39;
	13'hD5F: q=8'h7F;
	13'hD60: q=8'h0;
	13'hD61: q=8'h85;
	13'hD62: q=8'h37;
	13'hD63: q=8'h4F;
	13'hD64: q=8'hDD;
	13'hD65: q=8'h89;
	13'hD66: q=8'hDC;
	13'hD67: q=8'h9D;
	13'hD68: q=8'h93;
	13'hD69: q=8'h89;
	13'hD6A: q=8'h93;
	13'hD6B: q=8'h9B;
	13'hD6C: q=8'h25;
	13'hD6D: q=8'hB;
	13'hD6E: q=8'hD3;
	13'hD6F: q=8'h9B;
	13'hD70: q=8'hDD;
	13'hD71: q=8'h9D;
	13'hD72: q=8'hDE;
	13'hD73: q=8'h9D;
	13'hD74: q=8'h8;
	13'hD75: q=8'hDF;
	13'hD76: q=8'h9F;
	13'hD77: q=8'h33;
	13'hD78: q=8'h39;
	13'hD79: q=8'hC6;
	13'hD7A: q=8'h1A;
	13'hD7B: q=8'h73;
	13'hD7C: q=8'h0;
	13'hD7D: q=8'h85;
	13'hD7E: q=8'h27;
	13'hD7F: q=8'hC4;
	13'hD80: q=8'h8D;
	13'hD81: q=8'h3;
	13'hD82: q=8'h33;
	13'hD83: q=8'h20;
	13'hD84: q=8'hDD;
	13'hD85: q=8'hDE;
	13'hD86: q=8'hA1;
	13'hD87: q=8'hDF;
	13'hD88: q=8'h9D;
	13'hD89: q=8'h4F;
	13'hD8A: q=8'h5F;
	13'hD8B: q=8'hDD;
	13'hD8C: q=8'hC5;
	13'hD8D: q=8'hDE;
	13'hD8E: q=8'h9B;
	13'hD8F: q=8'hDF;
	13'hD90: q=8'hC1;
	13'hD91: q=8'hCE;
	13'hD92: q=8'h42;
	13'hD93: q=8'h41;
	13'hD94: q=8'hBC;
	13'hD95: q=8'h42;
	13'hD96: q=8'h3D;
	13'hD97: q=8'h27;
	13'hD98: q=8'h4;
	13'hD99: q=8'h8D;
	13'hD9A: q=8'h32;
	13'hD9B: q=8'h20;
	13'hD9C: q=8'hF7;
	13'hD9D: q=8'hDE;
	13'hD9E: q=8'h95;
	13'hD9F: q=8'h9C;
	13'hDA0: q=8'h97;
	13'hDA1: q=8'h27;
	13'hDA2: q=8'h4;
	13'hDA3: q=8'h8D;
	13'hDA4: q=8'h22;
	13'hDA5: q=8'h20;
	13'hDA6: q=8'hF8;
	13'hDA7: q=8'hDF;
	13'hDA8: q=8'hBB;
	13'hDA9: q=8'hDE;
	13'hDAA: q=8'hBB;
	13'hDAB: q=8'h9C;
	13'hDAC: q=8'h99;
	13'hDAD: q=8'h27;
	13'hDAE: q=8'h38;
	13'hDAF: q=8'hEC;
	13'hDB0: q=8'h2;
	13'hDB1: q=8'hD3;
	13'hDB2: q=8'hBB;
	13'hDB3: q=8'hDD;
	13'hDB4: q=8'hBB;
	13'hDB5: q=8'hA6;
	13'hDB6: q=8'h1;
	13'hDB7: q=8'h2A;
	13'hDB8: q=8'hF0;
	13'hDB9: q=8'hE6;
	13'hDBA: q=8'h4;
	13'hDBB: q=8'h58;
	13'hDBC: q=8'hCB;
	13'hDBD: q=8'h5;
	13'hDBE: q=8'h3A;
	13'hDBF: q=8'h9C;
	13'hDC0: q=8'hBB;
	13'hDC1: q=8'h27;
	13'hDC2: q=8'hE8;
	13'hDC3: q=8'h8D;
	13'hDC4: q=8'h8;
	13'hDC5: q=8'h20;
	13'hDC6: q=8'hF8;
	13'hDC7: q=8'hA6;
	13'hDC8: q=8'h1;
	13'hDC9: q=8'h8;
	13'hDCA: q=8'h8;
	13'hDCB: q=8'h2A;
	13'hDCC: q=8'h16;
	13'hDCD: q=8'hE6;
	13'hDCE: q=8'h0;
	13'hDCF: q=8'h27;
	13'hDD0: q=8'h12;
	13'hDD1: q=8'hEC;
	13'hDD2: q=8'h2;
	13'hDD3: q=8'h93;
	13'hDD4: q=8'h9D;
	13'hDD5: q=8'h22;
	13'hDD6: q=8'hC;
	13'hDD7: q=8'hEC;
	13'hDD8: q=8'h2;
	13'hDD9: q=8'h93;
	13'hDDA: q=8'hC1;
	13'hDDB: q=8'h23;
	13'hDDC: q=8'h6;
	13'hDDD: q=8'hDF;
	13'hDDE: q=8'hC5;
	13'hDDF: q=8'hEC;
	13'hDE0: q=8'h2;
	13'hDE1: q=8'hDD;
	13'hDE2: q=8'hC1;
	13'hDE3: q=8'hC6;
	13'hDE4: q=8'h5;
	13'hDE5: q=8'h3A;
	13'hDE6: q=8'h39;
	13'hDE7: q=8'hDE;
	13'hDE8: q=8'hC5;
	13'hDE9: q=8'h27;
	13'hDEA: q=8'hFB;
	13'hDEB: q=8'h4F;
	13'hDEC: q=8'hE6;
	13'hDED: q=8'h0;
	13'hDEE: q=8'h5A;
	13'hDEF: q=8'hD3;
	13'hDF0: q=8'hC1;
	13'hDF1: q=8'hDD;
	13'hDF2: q=8'hBD;
	13'hDF3: q=8'hDE;
	13'hDF4: q=8'h9D;
	13'hDF5: q=8'hDF;
	13'hDF6: q=8'hBB;
	13'hDF7: q=8'hBD;
	13'hDF8: q=8'hE2;
	13'hDF9: q=8'h0;
	13'hDFA: q=8'hDE;
	13'hDFB: q=8'hC5;
	13'hDFC: q=8'hDC;
	13'hDFD: q=8'hBF;
	13'hDFE: q=8'hED;
	13'hDFF: q=8'h2;
	13'hE00: q=8'hDE;
	13'hE01: q=8'hBF;
	13'hE02: q=8'h9;
	13'hE03: q=8'h7E;
	13'hE04: q=8'hED;
	13'hE05: q=8'h87;
	13'hE06: q=8'hDE;
	13'hE07: q=8'hCC;
	13'hE08: q=8'h3C;
	13'hE09: q=8'hBD;
	13'hE0A: q=8'hE9;
	13'hE0B: q=8'hE5;
	13'hE0C: q=8'hBD;
	13'hE0D: q=8'hE9;
	13'hE0E: q=8'hF;
	13'hE0F: q=8'h38;
	13'hE10: q=8'hDF;
	13'hE11: q=8'hDC;
	13'hE12: q=8'hE6;
	13'hE13: q=8'h0;
	13'hE14: q=8'hDE;
	13'hE15: q=8'hCC;
	13'hE16: q=8'hEB;
	13'hE17: q=8'h0;
	13'hE18: q=8'h24;
	13'hE19: q=8'h5;
	13'hE1A: q=8'hC6;
	13'hE1B: q=8'h1C;
	13'hE1C: q=8'h7E;
	13'hE1D: q=8'hE2;
	13'hE1E: q=8'h38;
	13'hE1F: q=8'hBD;
	13'hE20: q=8'hEC;
	13'hE21: q=8'hFC;
	13'hE22: q=8'hDE;
	13'hE23: q=8'hDC;
	13'hE24: q=8'hE6;
	13'hE25: q=8'h0;
	13'hE26: q=8'h8D;
	13'hE27: q=8'h10;
	13'hE28: q=8'hDE;
	13'hE29: q=8'hC7;
	13'hE2A: q=8'h8D;
	13'hE2B: q=8'h2C;
	13'hE2C: q=8'h8D;
	13'hE2D: q=8'hC;
	13'hE2E: q=8'hDE;
	13'hE2F: q=8'hDC;
	13'hE30: q=8'h8D;
	13'hE31: q=8'h26;
	13'hE32: q=8'hBD;
	13'hE33: q=8'hED;
	13'hE34: q=8'h3A;
	13'hE35: q=8'h7E;
	13'hE36: q=8'hE9;
	13'hE37: q=8'h2E;
	13'hE38: q=8'hEE;
	13'hE39: q=8'h2;
	13'hE3A: q=8'h7;
	13'hE3B: q=8'h36;
	13'hE3C: q=8'h9F;
	13'hE3D: q=8'h91;
	13'hE3E: q=8'hF;
	13'hE3F: q=8'h35;
	13'hE40: q=8'hDE;
	13'hE41: q=8'h9F;
	13'hE42: q=8'h5C;
	13'hE43: q=8'h20;
	13'hE44: q=8'h4;
	13'hE45: q=8'h32;
	13'hE46: q=8'hA7;
	13'hE47: q=8'h0;
	13'hE48: q=8'h8;
	13'hE49: q=8'h5A;
	13'hE4A: q=8'h26;
	13'hE4B: q=8'hF9;
	13'hE4C: q=8'hDF;
	13'hE4D: q=8'h9F;
	13'hE4E: q=8'h9E;
	13'hE4F: q=8'h91;
	13'hE50: q=8'h32;
	13'hE51: q=8'h6;
	13'hE52: q=8'h39;
	13'hE53: q=8'hBD;
	13'hE54: q=8'hE9;
	13'hE55: q=8'hF;
	13'hE56: q=8'hDE;
	13'hE57: q=8'hCC;
	13'hE58: q=8'hE6;
	13'hE59: q=8'h0;
	13'hE5A: q=8'h8D;
	13'hE5B: q=8'h14;
	13'hE5C: q=8'h26;
	13'hE5D: q=8'hF;
	13'hE5E: q=8'hEE;
	13'hE5F: q=8'h7;
	13'hE60: q=8'h9;
	13'hE61: q=8'h9C;
	13'hE62: q=8'h9D;
	13'hE63: q=8'h26;
	13'hE64: q=8'h6;
	13'hE65: q=8'h37;
	13'hE66: q=8'hD3;
	13'hE67: q=8'h9D;
	13'hE68: q=8'hDD;
	13'hE69: q=8'h9D;
	13'hE6A: q=8'h33;
	13'hE6B: q=8'h8;
	13'hE6C: q=8'h39;
	13'hE6D: q=8'hEE;
	13'hE6E: q=8'h2;
	13'hE6F: q=8'h39;
	13'hE70: q=8'hBC;
	13'hE71: q=8'h42;
	13'hE72: q=8'h3F;
	13'hE73: q=8'h26;
	13'hE74: q=8'hC;
	13'hE75: q=8'hFF;
	13'hE76: q=8'h42;
	13'hE77: q=8'h3D;
	13'hE78: q=8'h9;
	13'hE79: q=8'h9;
	13'hE7A: q=8'h9;
	13'hE7B: q=8'h9;
	13'hE7C: q=8'h9;
	13'hE7D: q=8'hFF;
	13'hE7E: q=8'h42;
	13'hE7F: q=8'h3F;
	13'hE80: q=8'h4F;
	13'hE81: q=8'h39;
	13'hE82: q=8'h8D;
	13'hE83: q=8'h3;
	13'hE84: q=8'h7E;
	13'hE85: q=8'hEC;
	13'hE86: q=8'hE2;
	13'hE87: q=8'h8D;
	13'hE88: q=8'hCA;
	13'hE89: q=8'h7F;
	13'hE8A: q=8'h0;
	13'hE8B: q=8'h84;
	13'hE8C: q=8'h5D;
	13'hE8D: q=8'h39;
	13'hE8E: q=8'hBD;
	13'hE8F: q=8'hEF;
	13'hE90: q=8'h10;
	13'hE91: q=8'hC6;
	13'hE92: q=8'h1;
	13'hE93: q=8'hBD;
	13'hE94: q=8'hED;
	13'hE95: q=8'h5F;
	13'hE96: q=8'h96;
	13'hE97: q=8'hCD;
	13'hE98: q=8'hBD;
	13'hE99: q=8'hED;
	13'hE9A: q=8'h0;
	13'hE9B: q=8'hA7;
	13'hE9C: q=8'h0;
	13'hE9D: q=8'h31;
	13'hE9E: q=8'h31;
	13'hE9F: q=8'h7E;
	13'hEA0: q=8'hED;
	13'hEA1: q=8'h3A;
	13'hEA2: q=8'h8D;
	13'hEA3: q=8'h2;
	13'hEA4: q=8'h20;
	13'hEA5: q=8'hDE;
	13'hEA6: q=8'h8D;
	13'hEA7: q=8'hDF;
	13'hEA8: q=8'h27;
	13'hEA9: q=8'h5D;
	13'hEAA: q=8'hE6;
	13'hEAB: q=8'h0;
	13'hEAC: q=8'h39;
	13'hEAD: q=8'h8D;
	13'hEAE: q=8'h43;
	13'hEAF: q=8'h4F;
	13'hEB0: q=8'hE1;
	13'hEB1: q=8'h0;
	13'hEB2: q=8'h23;
	13'hEB3: q=8'h3;
	13'hEB4: q=8'hE6;
	13'hEB5: q=8'h0;
	13'hEB6: q=8'h4F;
	13'hEB7: q=8'h37;
	13'hEB8: q=8'h36;
	13'hEB9: q=8'hBD;
	13'hEBA: q=8'hEC;
	13'hEBB: q=8'hFE;
	13'hEBC: q=8'hDE;
	13'hEBD: q=8'hC7;
	13'hEBE: q=8'h8D;
	13'hEBF: q=8'h98;
	13'hEC0: q=8'h33;
	13'hEC1: q=8'h3A;
	13'hEC2: q=8'h33;
	13'hEC3: q=8'hBD;
	13'hEC4: q=8'hEE;
	13'hEC5: q=8'h3A;
	13'hEC6: q=8'h20;
	13'hEC7: q=8'hD7;
	13'hEC8: q=8'h8D;
	13'hEC9: q=8'h28;
	13'hECA: q=8'hA6;
	13'hECB: q=8'h0;
	13'hECC: q=8'h10;
	13'hECD: q=8'h20;
	13'hECE: q=8'hE1;
	13'hECF: q=8'hC6;
	13'hED0: q=8'hFF;
	13'hED1: q=8'hD7;
	13'hED2: q=8'hCD;
	13'hED3: q=8'h8D;
	13'hED4: q=8'h44;
	13'hED5: q=8'h81;
	13'hED6: q=8'h29;
	13'hED7: q=8'h27;
	13'hED8: q=8'h3;
	13'hED9: q=8'hBD;
	13'hEDA: q=8'hEF;
	13'hEDB: q=8'h47;
	13'hEDC: q=8'h8D;
	13'hEDD: q=8'h14;
	13'hEDE: q=8'h27;
	13'hEDF: q=8'h27;
	13'hEE0: q=8'h5F;
	13'hEE1: q=8'h4A;
	13'hEE2: q=8'hA1;
	13'hEE3: q=8'h0;
	13'hEE4: q=8'h24;
	13'hEE5: q=8'hD1;
	13'hEE6: q=8'h16;
	13'hEE7: q=8'hE0;
	13'hEE8: q=8'h0;
	13'hEE9: q=8'h50;
	13'hEEA: q=8'hD1;
	13'hEEB: q=8'hCD;
	13'hEEC: q=8'h23;
	13'hEED: q=8'hC9;
	13'hEEE: q=8'hD6;
	13'hEEF: q=8'hCD;
	13'hEF0: q=8'h20;
	13'hEF1: q=8'hC5;
	13'hEF2: q=8'hBD;
	13'hEF3: q=8'hEA;
	13'hEF4: q=8'h29;
	13'hEF5: q=8'h30;
	13'hEF6: q=8'hEC;
	13'hEF7: q=8'h5;
	13'hEF8: q=8'hDD;
	13'hEF9: q=8'hC7;
	13'hEFA: q=8'hEC;
	13'hEFB: q=8'h0;
	13'hEFC: q=8'hED;
	13'hEFD: q=8'h5;
	13'hEFE: q=8'h31;
	13'hEFF: q=8'h31;
	13'hF00: q=8'h31;
	13'hF01: q=8'h31;
	13'hF02: q=8'h32;
	13'hF03: q=8'hDE;
	13'hF04: q=8'hC7;
	13'hF05: q=8'h16;
	13'hF06: q=8'h39;
	13'hF07: q=8'h7E;
	13'hF08: q=8'hEC;
	13'hF09: q=8'h2E;
	13'hF0A: q=8'hBD;
	13'hF0B: q=8'h0;
	13'hF0C: q=8'hEB;
	13'hF0D: q=8'hBD;
	13'hF0E: q=8'hE9;
	13'hF0F: q=8'hC;
	13'hF10: q=8'hBD;
	13'hF11: q=8'hEB;
	13'hF12: q=8'hC0;
	13'hF13: q=8'h96;
	13'hF14: q=8'hCC;
	13'hF15: q=8'h26;
	13'hF16: q=8'hF0;
	13'hF17: q=8'hD6;
	13'hF18: q=8'hCD;
	13'hF19: q=8'h7E;
	13'hF1A: q=8'h0;
	13'hF1B: q=8'hF3;
	13'hF1C: q=8'hBD;
	13'hF1D: q=8'hEE;
	13'hF1E: q=8'h87;
	13'hF1F: q=8'h26;
	13'hF20: q=8'h3;
	13'hF21: q=8'h7E;
	13'hF22: q=8'hEF;
	13'hF23: q=8'hF4;
	13'hF24: q=8'hBD;
	13'hF25: q=8'hE2;
	13'hF26: q=8'h2C;
	13'hF27: q=8'hA6;
	13'hF28: q=8'h0;
	13'hF29: q=8'h36;
	13'hF2A: q=8'h6F;
	13'hF2B: q=8'h0;
	13'hF2C: q=8'hDE;
	13'hF2D: q=8'hF4;
	13'hF2E: q=8'hDF;
	13'hF2F: q=8'hDE;
	13'hF30: q=8'hDE;
	13'hF31: q=8'h89;
	13'hF32: q=8'hDF;
	13'hF33: q=8'hF4;
	13'hF34: q=8'h8D;
	13'hF35: q=8'hE3;
	13'hF36: q=8'hBD;
	13'hF37: q=8'hF3;
	13'hF38: q=8'h59;
	13'hF39: q=8'h32;
	13'hF3A: q=8'hDE;
	13'hF3B: q=8'h8B;
	13'hF3C: q=8'hA7;
	13'hF3D: q=8'h0;
	13'hF3E: q=8'hDE;
	13'hF3F: q=8'hDE;
	13'hF40: q=8'hDF;
	13'hF41: q=8'hF4;
	13'hF42: q=8'h39;
	13'hF43: q=8'h8D;
	13'hF44: q=8'h7;
	13'hF45: q=8'hDF;
	13'hF46: q=8'hA5;
	13'hF47: q=8'hBD;
	13'hF48: q=8'hEA;
	13'hF49: q=8'h2F;
	13'hF4A: q=8'h20;
	13'hF4B: q=8'hC1;
	13'hF4C: q=8'hBD;
	13'hF4D: q=8'hE9;
	13'hF4E: q=8'hC;
	13'hF4F: q=8'h96;
	13'hF50: q=8'hCE;
	13'hF51: q=8'h2B;
	13'hF52: q=8'hB4;
	13'hF53: q=8'h96;
	13'hF54: q=8'hC9;
	13'hF55: q=8'h81;
	13'hF56: q=8'h90;
	13'hF57: q=8'h22;
	13'hF58: q=8'hAE;
	13'hF59: q=8'hBD;
	13'hF5A: q=8'hF3;
	13'hF5B: q=8'hB;
	13'hF5C: q=8'hDE;
	13'hF5D: q=8'hCC;
	13'hF5E: q=8'h39;
	13'hF5F: q=8'h8D;
	13'hF60: q=8'hEE;
	13'hF61: q=8'hE6;
	13'hF62: q=8'h0;
	13'hF63: q=8'h7E;
	13'hF64: q=8'hEC;
	13'hF65: q=8'hE2;
	13'hF66: q=8'h8D;
	13'hF67: q=8'hDB;
	13'hF68: q=8'hDE;
	13'hF69: q=8'hA5;
	13'hF6A: q=8'hE7;
	13'hF6B: q=8'h0;
	13'hF6C: q=8'h39;
	13'hF6D: q=8'hCE;
	13'hF6E: q=8'hF5;
	13'hF6F: q=8'h24;
	13'hF70: q=8'h20;
	13'hF71: q=8'hB;
	13'hF72: q=8'hBD;
	13'hF73: q=8'hF1;
	13'hF74: q=8'h60;
	13'hF75: q=8'h73;
	13'hF76: q=8'h0;
	13'hF77: q=8'hCE;
	13'hF78: q=8'h73;
	13'hF79: q=8'h0;
	13'hF7A: q=8'hDC;
	13'hF7B: q=8'h20;
	13'hF7C: q=8'h3;
	13'hF7D: q=8'hBD;
	13'hF7E: q=8'hF1;
	13'hF7F: q=8'h60;
	13'hF80: q=8'h5D;
	13'hF81: q=8'h26;
	13'hF82: q=8'h3;
	13'hF83: q=8'h7E;
	13'hF84: q=8'hF2;
	13'hF85: q=8'h8B;
	13'hF86: q=8'hCE;
	13'hF87: q=8'h0;
	13'hF88: q=8'hD6;
	13'hF89: q=8'h16;
	13'hF8A: q=8'h27;
	13'hF8B: q=8'h6D;
	13'hF8C: q=8'hD0;
	13'hF8D: q=8'hC9;
	13'hF8E: q=8'h27;
	13'hF8F: q=8'h6A;
	13'hF90: q=8'h2B;
	13'hF91: q=8'hA;
	13'hF92: q=8'h97;
	13'hF93: q=8'hC9;
	13'hF94: q=8'h96;
	13'hF95: q=8'hDB;
	13'hF96: q=8'h97;
	13'hF97: q=8'hCE;
	13'hF98: q=8'hCE;
	13'hF99: q=8'h0;
	13'hF9A: q=8'hC9;
	13'hF9B: q=8'h50;
	13'hF9C: q=8'hC1;
	13'hF9D: q=8'hF8;
	13'hF9E: q=8'h2F;
	13'hF9F: q=8'h5A;
	13'hFA0: q=8'h4F;
	13'hFA1: q=8'h64;
	13'hFA2: q=8'h1;
	13'hFA3: q=8'hBD;
	13'hFA4: q=8'hF0;
	13'hFA5: q=8'h80;
	13'hFA6: q=8'hD6;
	13'hFA7: q=8'hDC;
	13'hFA8: q=8'h2A;
	13'hFA9: q=8'hB;
	13'hFAA: q=8'h63;
	13'hFAB: q=8'h1;
	13'hFAC: q=8'h63;
	13'hFAD: q=8'h2;
	13'hFAE: q=8'h63;
	13'hFAF: q=8'h3;
	13'hFB0: q=8'h63;
	13'hFB1: q=8'h4;
	13'hFB2: q=8'h43;
	13'hFB3: q=8'h89;
	13'hFB4: q=8'h0;
	13'hFB5: q=8'h97;
	13'hFB6: q=8'hDD;
	13'hFB7: q=8'h96;
	13'hFB8: q=8'hCD;
	13'hFB9: q=8'h99;
	13'hFBA: q=8'hDA;
	13'hFBB: q=8'h97;
	13'hFBC: q=8'hCD;
	13'hFBD: q=8'h96;
	13'hFBE: q=8'hCC;
	13'hFBF: q=8'h99;
	13'hFC0: q=8'hD9;
	13'hFC1: q=8'h97;
	13'hFC2: q=8'hCC;
	13'hFC3: q=8'h96;
	13'hFC4: q=8'hCB;
	13'hFC5: q=8'h99;
	13'hFC6: q=8'hD8;
	13'hFC7: q=8'h97;
	13'hFC8: q=8'hCB;
	13'hFC9: q=8'h96;
	13'hFCA: q=8'hCA;
	13'hFCB: q=8'h99;
	13'hFCC: q=8'hD7;
	13'hFCD: q=8'h97;
	13'hFCE: q=8'hCA;
	13'hFCF: q=8'h17;
	13'hFD0: q=8'h2A;
	13'hFD1: q=8'h47;
	13'hFD2: q=8'h25;
	13'hFD3: q=8'h2;
	13'hFD4: q=8'h8D;
	13'hFD5: q=8'h66;
	13'hFD6: q=8'h5F;
	13'hFD7: q=8'h96;
	13'hFD8: q=8'hCA;
	13'hFD9: q=8'h26;
	13'hFDA: q=8'h34;
	13'hFDB: q=8'h96;
	13'hFDC: q=8'hCB;
	13'hFDD: q=8'h97;
	13'hFDE: q=8'hCA;
	13'hFDF: q=8'h96;
	13'hFE0: q=8'hCC;
	13'hFE1: q=8'h97;
	13'hFE2: q=8'hCB;
	13'hFE3: q=8'h96;
	13'hFE4: q=8'hCD;
	13'hFE5: q=8'h97;
	13'hFE6: q=8'hCC;
	13'hFE7: q=8'h96;
	13'hFE8: q=8'hDD;
	13'hFE9: q=8'h97;
	13'hFEA: q=8'hCD;
	13'hFEB: q=8'h7F;
	13'hFEC: q=8'h0;
	13'hFED: q=8'hDD;
	13'hFEE: q=8'hCB;
	13'hFEF: q=8'h8;
	13'hFF0: q=8'hC1;
	13'hFF1: q=8'h28;
	13'hFF2: q=8'h2D;
	13'hFF3: q=8'hE3;
	13'hFF4: q=8'h4F;
	13'hFF5: q=8'h97;
	13'hFF6: q=8'hC9;
	13'hFF7: q=8'h97;
	13'hFF8: q=8'hCE;
	13'hFF9: q=8'h39;
	13'hFFA: q=8'h8D;
	13'hFFB: q=8'h78;
	13'hFFC: q=8'hC;
	13'hFFD: q=8'h20;
	13'hFFE: q=8'hA7;
	13'hFFF: q=8'h5C;
	13'h1000: q=8'h78;
	13'h1001: q=8'h0;
	13'h1002: q=8'hDD;
	13'h1003: q=8'h79;
	13'h1004: q=8'h0;
	13'h1005: q=8'hCD;
	13'h1006: q=8'h79;
	13'h1007: q=8'h0;
	13'h1008: q=8'hCC;
	13'h1009: q=8'h79;
	13'h100A: q=8'h0;
	13'h100B: q=8'hCB;
	13'h100C: q=8'h79;
	13'h100D: q=8'h0;
	13'h100E: q=8'hCA;
	13'h100F: q=8'h2A;
	13'h1010: q=8'hEE;
	13'h1011: q=8'h96;
	13'h1012: q=8'hC9;
	13'h1013: q=8'h10;
	13'h1014: q=8'h97;
	13'h1015: q=8'hC9;
	13'h1016: q=8'h23;
	13'h1017: q=8'hDC;
	13'h1018: q=8'h8C;
	13'h1019: q=8'h25;
	13'h101A: q=8'h9;
	13'h101B: q=8'h78;
	13'h101C: q=8'h0;
	13'h101D: q=8'hDD;
	13'h101E: q=8'h86;
	13'h101F: q=8'h0;
	13'h1020: q=8'h97;
	13'h1021: q=8'hDD;
	13'h1022: q=8'h20;
	13'h1023: q=8'h11;
	13'h1024: q=8'h7C;
	13'h1025: q=8'h0;
	13'h1026: q=8'hC9;
	13'h1027: q=8'h27;
	13'h1028: q=8'h2F;
	13'h1029: q=8'h76;
	13'h102A: q=8'h0;
	13'h102B: q=8'hCA;
	13'h102C: q=8'h76;
	13'h102D: q=8'h0;
	13'h102E: q=8'hCB;
	13'h102F: q=8'h76;
	13'h1030: q=8'h0;
	13'h1031: q=8'hCC;
	13'h1032: q=8'h76;
	13'h1033: q=8'h0;
	13'h1034: q=8'hCD;
	13'h1035: q=8'h24;
	13'h1036: q=8'h4;
	13'h1037: q=8'h8D;
	13'h1038: q=8'h12;
	13'h1039: q=8'h27;
	13'h103A: q=8'hE9;
	13'h103B: q=8'h39;
	13'h103C: q=8'h73;
	13'h103D: q=8'h0;
	13'h103E: q=8'hCE;
	13'h103F: q=8'h73;
	13'h1040: q=8'h0;
	13'h1041: q=8'hCA;
	13'h1042: q=8'h73;
	13'h1043: q=8'h0;
	13'h1044: q=8'hCB;
	13'h1045: q=8'h73;
	13'h1046: q=8'h0;
	13'h1047: q=8'hCC;
	13'h1048: q=8'h73;
	13'h1049: q=8'h0;
	13'h104A: q=8'hCD;
	13'h104B: q=8'hDE;
	13'h104C: q=8'hCC;
	13'h104D: q=8'h8;
	13'h104E: q=8'hDF;
	13'h104F: q=8'hCC;
	13'h1050: q=8'h26;
	13'h1051: q=8'h5;
	13'h1052: q=8'hDE;
	13'h1053: q=8'hCA;
	13'h1054: q=8'h8;
	13'h1055: q=8'hDF;
	13'h1056: q=8'hCA;
	13'h1057: q=8'h39;
	13'h1058: q=8'hC6;
	13'h1059: q=8'hA;
	13'h105A: q=8'h7E;
	13'h105B: q=8'hE2;
	13'h105C: q=8'h38;
	13'h105D: q=8'hCE;
	13'h105E: q=8'h0;
	13'h105F: q=8'h8C;
	13'h1060: q=8'hA6;
	13'h1061: q=8'h4;
	13'h1062: q=8'h97;
	13'h1063: q=8'hDD;
	13'h1064: q=8'hA6;
	13'h1065: q=8'h3;
	13'h1066: q=8'hA7;
	13'h1067: q=8'h4;
	13'h1068: q=8'hA6;
	13'h1069: q=8'h2;
	13'h106A: q=8'hA7;
	13'h106B: q=8'h3;
	13'h106C: q=8'hA6;
	13'h106D: q=8'h1;
	13'h106E: q=8'hA7;
	13'h106F: q=8'h2;
	13'h1070: q=8'h96;
	13'h1071: q=8'hD5;
	13'h1072: q=8'hA7;
	13'h1073: q=8'h1;
	13'h1074: q=8'hCB;
	13'h1075: q=8'h8;
	13'h1076: q=8'h2F;
	13'h1077: q=8'hE8;
	13'h1078: q=8'h96;
	13'h1079: q=8'hDD;
	13'h107A: q=8'hC0;
	13'h107B: q=8'h8;
	13'h107C: q=8'h27;
	13'h107D: q=8'hC;
	13'h107E: q=8'h67;
	13'h107F: q=8'h1;
	13'h1080: q=8'h66;
	13'h1081: q=8'h2;
	13'h1082: q=8'h66;
	13'h1083: q=8'h3;
	13'h1084: q=8'h66;
	13'h1085: q=8'h4;
	13'h1086: q=8'h46;
	13'h1087: q=8'h5C;
	13'h1088: q=8'h26;
	13'h1089: q=8'hF4;
	13'h108A: q=8'h39;
	13'h108B: q=8'h81;
	13'h108C: q=8'h0;
	13'h108D: q=8'h0;
	13'h108E: q=8'h0;
	13'h108F: q=8'h0;
	13'h1090: q=8'h3;
	13'h1091: q=8'h7F;
	13'h1092: q=8'h5E;
	13'h1093: q=8'h56;
	13'h1094: q=8'hCB;
	13'h1095: q=8'h79;
	13'h1096: q=8'h80;
	13'h1097: q=8'h13;
	13'h1098: q=8'h9B;
	13'h1099: q=8'hB;
	13'h109A: q=8'h64;
	13'h109B: q=8'h80;
	13'h109C: q=8'h76;
	13'h109D: q=8'h38;
	13'h109E: q=8'h93;
	13'h109F: q=8'h16;
	13'h10A0: q=8'h82;
	13'h10A1: q=8'h38;
	13'h10A2: q=8'hAA;
	13'h10A3: q=8'h3B;
	13'h10A4: q=8'h20;
	13'h10A5: q=8'h80;
	13'h10A6: q=8'h35;
	13'h10A7: q=8'h4;
	13'h10A8: q=8'hF3;
	13'h10A9: q=8'h34;
	13'h10AA: q=8'h81;
	13'h10AB: q=8'h35;
	13'h10AC: q=8'h4;
	13'h10AD: q=8'hF3;
	13'h10AE: q=8'h34;
	13'h10AF: q=8'h80;
	13'h10B0: q=8'h80;
	13'h10B1: q=8'h0;
	13'h10B2: q=8'h0;
	13'h10B3: q=8'h0;
	13'h10B4: q=8'h80;
	13'h10B5: q=8'h31;
	13'h10B6: q=8'h72;
	13'h10B7: q=8'h17;
	13'h10B8: q=8'hF8;
	13'h10B9: q=8'hBD;
	13'h10BA: q=8'hF2;
	13'h10BB: q=8'hAD;
	13'h10BC: q=8'h2E;
	13'h10BD: q=8'h3;
	13'h10BE: q=8'h7E;
	13'h10BF: q=8'hEC;
	13'h10C0: q=8'h2E;
	13'h10C1: q=8'hCE;
	13'h10C2: q=8'hF0;
	13'h10C3: q=8'hA5;
	13'h10C4: q=8'h96;
	13'h10C5: q=8'hC9;
	13'h10C6: q=8'h80;
	13'h10C7: q=8'h80;
	13'h10C8: q=8'h36;
	13'h10C9: q=8'h86;
	13'h10CA: q=8'h80;
	13'h10CB: q=8'h97;
	13'h10CC: q=8'hC9;
	13'h10CD: q=8'hBD;
	13'h10CE: q=8'hEF;
	13'h10CF: q=8'h7D;
	13'h10D0: q=8'hCE;
	13'h10D1: q=8'hF0;
	13'h10D2: q=8'hAA;
	13'h10D3: q=8'hBD;
	13'h10D4: q=8'hF1;
	13'h10D5: q=8'hC6;
	13'h10D6: q=8'hCE;
	13'h10D7: q=8'hF0;
	13'h10D8: q=8'h8B;
	13'h10D9: q=8'hBD;
	13'h10DA: q=8'hEF;
	13'h10DB: q=8'h72;
	13'h10DC: q=8'hCE;
	13'h10DD: q=8'hF0;
	13'h10DE: q=8'h90;
	13'h10DF: q=8'hBD;
	13'h10E0: q=8'hF5;
	13'h10E1: q=8'hF8;
	13'h10E2: q=8'hCE;
	13'h10E3: q=8'hF0;
	13'h10E4: q=8'hAF;
	13'h10E5: q=8'hBD;
	13'h10E6: q=8'hEF;
	13'h10E7: q=8'h7D;
	13'h10E8: q=8'h33;
	13'h10E9: q=8'hBD;
	13'h10EA: q=8'hF3;
	13'h10EB: q=8'hE9;
	13'h10EC: q=8'hCE;
	13'h10ED: q=8'hF0;
	13'h10EE: q=8'hB4;
	13'h10EF: q=8'h8D;
	13'h10F0: q=8'h6F;
	13'h10F1: q=8'h27;
	13'h10F2: q=8'h6C;
	13'h10F3: q=8'hBD;
	13'h10F4: q=8'hF1;
	13'h10F5: q=8'h79;
	13'h10F6: q=8'h86;
	13'h10F7: q=8'h0;
	13'h10F8: q=8'h97;
	13'h10F9: q=8'h8D;
	13'h10FA: q=8'h97;
	13'h10FB: q=8'h8E;
	13'h10FC: q=8'h97;
	13'h10FD: q=8'h8F;
	13'h10FE: q=8'h97;
	13'h10FF: q=8'h90;
	13'h1100: q=8'hD6;
	13'h1101: q=8'hCD;
	13'h1102: q=8'h8D;
	13'h1103: q=8'h26;
	13'h1104: q=8'hD6;
	13'h1105: q=8'hDD;
	13'h1106: q=8'hF7;
	13'h1107: q=8'h42;
	13'h1108: q=8'h55;
	13'h1109: q=8'hD6;
	13'h110A: q=8'hCC;
	13'h110B: q=8'h8D;
	13'h110C: q=8'h1D;
	13'h110D: q=8'hD6;
	13'h110E: q=8'hDD;
	13'h110F: q=8'hF7;
	13'h1110: q=8'h42;
	13'h1111: q=8'h54;
	13'h1112: q=8'hD6;
	13'h1113: q=8'hCB;
	13'h1114: q=8'h8D;
	13'h1115: q=8'h14;
	13'h1116: q=8'hD6;
	13'h1117: q=8'hDD;
	13'h1118: q=8'hF7;
	13'h1119: q=8'h42;
	13'h111A: q=8'h53;
	13'h111B: q=8'hD6;
	13'h111C: q=8'hCA;
	13'h111D: q=8'h8D;
	13'h111E: q=8'h10;
	13'h111F: q=8'hD6;
	13'h1120: q=8'hDD;
	13'h1121: q=8'hF7;
	13'h1122: q=8'h42;
	13'h1123: q=8'h52;
	13'h1124: q=8'hBD;
	13'h1125: q=8'hF2;
	13'h1126: q=8'h48;
	13'h1127: q=8'h7E;
	13'h1128: q=8'hEF;
	13'h1129: q=8'hD6;
	13'h112A: q=8'h26;
	13'h112B: q=8'h3;
	13'h112C: q=8'h7E;
	13'h112D: q=8'hF0;
	13'h112E: q=8'h5D;
	13'h112F: q=8'hD;
	13'h1130: q=8'h96;
	13'h1131: q=8'h8D;
	13'h1132: q=8'h56;
	13'h1133: q=8'h27;
	13'h1134: q=8'h2A;
	13'h1135: q=8'h24;
	13'h1136: q=8'h16;
	13'h1137: q=8'h96;
	13'h1138: q=8'h90;
	13'h1139: q=8'h9B;
	13'h113A: q=8'hDA;
	13'h113B: q=8'h97;
	13'h113C: q=8'h90;
	13'h113D: q=8'h96;
	13'h113E: q=8'h8F;
	13'h113F: q=8'h99;
	13'h1140: q=8'hD9;
	13'h1141: q=8'h97;
	13'h1142: q=8'h8F;
	13'h1143: q=8'h96;
	13'h1144: q=8'h8E;
	13'h1145: q=8'h99;
	13'h1146: q=8'hD8;
	13'h1147: q=8'h97;
	13'h1148: q=8'h8E;
	13'h1149: q=8'h96;
	13'h114A: q=8'h8D;
	13'h114B: q=8'h99;
	13'h114C: q=8'hD7;
	13'h114D: q=8'h46;
	13'h114E: q=8'h97;
	13'h114F: q=8'h8D;
	13'h1150: q=8'h76;
	13'h1151: q=8'h0;
	13'h1152: q=8'h8E;
	13'h1153: q=8'h76;
	13'h1154: q=8'h0;
	13'h1155: q=8'h8F;
	13'h1156: q=8'h76;
	13'h1157: q=8'h0;
	13'h1158: q=8'h90;
	13'h1159: q=8'h76;
	13'h115A: q=8'h0;
	13'h115B: q=8'hDD;
	13'h115C: q=8'hC;
	13'h115D: q=8'h20;
	13'h115E: q=8'hD1;
	13'h115F: q=8'h39;
	13'h1160: q=8'hEC;
	13'h1161: q=8'h1;
	13'h1162: q=8'h97;
	13'h1163: q=8'hDB;
	13'h1164: q=8'h8A;
	13'h1165: q=8'h80;
	13'h1166: q=8'hDD;
	13'h1167: q=8'hD7;
	13'h1168: q=8'hD6;
	13'h1169: q=8'hDB;
	13'h116A: q=8'hD8;
	13'h116B: q=8'hCE;
	13'h116C: q=8'hD7;
	13'h116D: q=8'hDC;
	13'h116E: q=8'hEC;
	13'h116F: q=8'h3;
	13'h1170: q=8'hDD;
	13'h1171: q=8'hD9;
	13'h1172: q=8'hA6;
	13'h1173: q=8'h0;
	13'h1174: q=8'h97;
	13'h1175: q=8'hD6;
	13'h1176: q=8'hD6;
	13'h1177: q=8'hC9;
	13'h1178: q=8'h39;
	13'h1179: q=8'h4D;
	13'h117A: q=8'h27;
	13'h117B: q=8'h19;
	13'h117C: q=8'h9B;
	13'h117D: q=8'hC9;
	13'h117E: q=8'h46;
	13'h117F: q=8'h49;
	13'h1180: q=8'h28;
	13'h1181: q=8'h13;
	13'h1182: q=8'h8B;
	13'h1183: q=8'h80;
	13'h1184: q=8'h97;
	13'h1185: q=8'hC9;
	13'h1186: q=8'h26;
	13'h1187: q=8'h3;
	13'h1188: q=8'h7E;
	13'h1189: q=8'hEF;
	13'h118A: q=8'hF7;
	13'h118B: q=8'h96;
	13'h118C: q=8'hDC;
	13'h118D: q=8'h97;
	13'h118E: q=8'hCE;
	13'h118F: q=8'h39;
	13'h1190: q=8'h96;
	13'h1191: q=8'hCE;
	13'h1192: q=8'h43;
	13'h1193: q=8'h20;
	13'h1194: q=8'h2;
	13'h1195: q=8'h32;
	13'h1196: q=8'h32;
	13'h1197: q=8'h2B;
	13'h1198: q=8'h3;
	13'h1199: q=8'h7E;
	13'h119A: q=8'hEF;
	13'h119B: q=8'hF4;
	13'h119C: q=8'h7E;
	13'h119D: q=8'hF0;
	13'h119E: q=8'h58;
	13'h119F: q=8'hBD;
	13'h11A0: q=8'hF2;
	13'h11A1: q=8'h9F;
	13'h11A2: q=8'h27;
	13'h11A3: q=8'hF;
	13'h11A4: q=8'h8B;
	13'h11A5: q=8'h2;
	13'h11A6: q=8'h25;
	13'h11A7: q=8'hF4;
	13'h11A8: q=8'h7F;
	13'h11A9: q=8'h0;
	13'h11AA: q=8'hDC;
	13'h11AB: q=8'hBD;
	13'h11AC: q=8'hEF;
	13'h11AD: q=8'h89;
	13'h11AE: q=8'h7C;
	13'h11AF: q=8'h0;
	13'h11B0: q=8'hC9;
	13'h11B1: q=8'h27;
	13'h11B2: q=8'hE9;
	13'h11B3: q=8'h39;
	13'h11B4: q=8'h84;
	13'h11B5: q=8'h20;
	13'h11B6: q=8'h0;
	13'h11B7: q=8'h0;
	13'h11B8: q=8'h0;
	13'h11B9: q=8'hBD;
	13'h11BA: q=8'hF2;
	13'h11BB: q=8'h9F;
	13'h11BC: q=8'hCE;
	13'h11BD: q=8'hF1;
	13'h11BE: q=8'hB4;
	13'h11BF: q=8'h5F;
	13'h11C0: q=8'hD7;
	13'h11C1: q=8'hDC;
	13'h11C2: q=8'hBD;
	13'h11C3: q=8'hF2;
	13'h11C4: q=8'h51;
	13'h11C5: q=8'h8C;
	13'h11C6: q=8'h8D;
	13'h11C7: q=8'h98;
	13'h11C8: q=8'h27;
	13'h11C9: q=8'h79;
	13'h11CA: q=8'h70;
	13'h11CB: q=8'h0;
	13'h11CC: q=8'hC9;
	13'h11CD: q=8'h8D;
	13'h11CE: q=8'hAA;
	13'h11CF: q=8'h7C;
	13'h11D0: q=8'h0;
	13'h11D1: q=8'hC9;
	13'h11D2: q=8'h27;
	13'h11D3: q=8'hC8;
	13'h11D4: q=8'hCE;
	13'h11D5: q=8'h0;
	13'h11D6: q=8'h8D;
	13'h11D7: q=8'hC6;
	13'h11D8: q=8'h4;
	13'h11D9: q=8'hD7;
	13'h11DA: q=8'h82;
	13'h11DB: q=8'hC6;
	13'h11DC: q=8'h1;
	13'h11DD: q=8'h96;
	13'h11DE: q=8'hCA;
	13'h11DF: q=8'h91;
	13'h11E0: q=8'hD7;
	13'h11E1: q=8'h26;
	13'h11E2: q=8'h13;
	13'h11E3: q=8'h96;
	13'h11E4: q=8'hCB;
	13'h11E5: q=8'h91;
	13'h11E6: q=8'hD8;
	13'h11E7: q=8'h26;
	13'h11E8: q=8'hD;
	13'h11E9: q=8'h96;
	13'h11EA: q=8'hCC;
	13'h11EB: q=8'h91;
	13'h11EC: q=8'hD9;
	13'h11ED: q=8'h26;
	13'h11EE: q=8'h7;
	13'h11EF: q=8'h96;
	13'h11F0: q=8'hCD;
	13'h11F1: q=8'h91;
	13'h11F2: q=8'hDA;
	13'h11F3: q=8'h26;
	13'h11F4: q=8'h1;
	13'h11F5: q=8'hD;
	13'h11F6: q=8'h7;
	13'h11F7: q=8'h59;
	13'h11F8: q=8'h24;
	13'h11F9: q=8'hC;
	13'h11FA: q=8'hE7;
	13'h11FB: q=8'h0;
	13'h11FC: q=8'h8;
	13'h11FD: q=8'h7A;
	13'h11FE: q=8'h0;
	13'h11FF: q=8'h82;
	13'h1200: q=8'h2B;
	13'h1201: q=8'h37;
	13'h1202: q=8'h27;
	13'h1203: q=8'h31;
	13'h1204: q=8'hC6;
	13'h1205: q=8'h1;
	13'h1206: q=8'h6;
	13'h1207: q=8'h25;
	13'h1208: q=8'h12;
	13'h1209: q=8'h78;
	13'h120A: q=8'h0;
	13'h120B: q=8'hDA;
	13'h120C: q=8'h79;
	13'h120D: q=8'h0;
	13'h120E: q=8'hD9;
	13'h120F: q=8'h79;
	13'h1210: q=8'h0;
	13'h1211: q=8'hD8;
	13'h1212: q=8'h79;
	13'h1213: q=8'h0;
	13'h1214: q=8'hD7;
	13'h1215: q=8'h25;
	13'h1216: q=8'hDF;
	13'h1217: q=8'h2B;
	13'h1218: q=8'hC4;
	13'h1219: q=8'h20;
	13'h121A: q=8'hDB;
	13'h121B: q=8'h96;
	13'h121C: q=8'hDA;
	13'h121D: q=8'h90;
	13'h121E: q=8'hCD;
	13'h121F: q=8'h97;
	13'h1220: q=8'hDA;
	13'h1221: q=8'h96;
	13'h1222: q=8'hD9;
	13'h1223: q=8'h92;
	13'h1224: q=8'hCC;
	13'h1225: q=8'h97;
	13'h1226: q=8'hD9;
	13'h1227: q=8'h96;
	13'h1228: q=8'hD8;
	13'h1229: q=8'h92;
	13'h122A: q=8'hCB;
	13'h122B: q=8'h97;
	13'h122C: q=8'hD8;
	13'h122D: q=8'h96;
	13'h122E: q=8'hD7;
	13'h122F: q=8'h92;
	13'h1230: q=8'hCA;
	13'h1231: q=8'h97;
	13'h1232: q=8'hD7;
	13'h1233: q=8'h20;
	13'h1234: q=8'hD4;
	13'h1235: q=8'hC6;
	13'h1236: q=8'h40;
	13'h1237: q=8'h20;
	13'h1238: q=8'hCD;
	13'h1239: q=8'h56;
	13'h123A: q=8'h56;
	13'h123B: q=8'h56;
	13'h123C: q=8'hD7;
	13'h123D: q=8'hDD;
	13'h123E: q=8'h8D;
	13'h123F: q=8'h8;
	13'h1240: q=8'h7E;
	13'h1241: q=8'hEF;
	13'h1242: q=8'hD6;
	13'h1243: q=8'hC6;
	13'h1244: q=8'h14;
	13'h1245: q=8'h7E;
	13'h1246: q=8'hE2;
	13'h1247: q=8'h38;
	13'h1248: q=8'hDE;
	13'h1249: q=8'h8D;
	13'h124A: q=8'hDF;
	13'h124B: q=8'hCA;
	13'h124C: q=8'hDE;
	13'h124D: q=8'h8F;
	13'h124E: q=8'hDF;
	13'h124F: q=8'hCC;
	13'h1250: q=8'h39;
	13'h1251: q=8'h36;
	13'h1252: q=8'hEC;
	13'h1253: q=8'h1;
	13'h1254: q=8'h97;
	13'h1255: q=8'hCE;
	13'h1256: q=8'h8A;
	13'h1257: q=8'h80;
	13'h1258: q=8'hDD;
	13'h1259: q=8'hCA;
	13'h125A: q=8'h7F;
	13'h125B: q=8'h0;
	13'h125C: q=8'hDD;
	13'h125D: q=8'hE6;
	13'h125E: q=8'h0;
	13'h125F: q=8'hEE;
	13'h1260: q=8'h3;
	13'h1261: q=8'hDF;
	13'h1262: q=8'hCC;
	13'h1263: q=8'hD7;
	13'h1264: q=8'hC9;
	13'h1265: q=8'h32;
	13'h1266: q=8'h39;
	13'h1267: q=8'hCE;
	13'h1268: q=8'h0;
	13'h1269: q=8'hBF;
	13'h126A: q=8'h20;
	13'h126B: q=8'h6;
	13'h126C: q=8'hCE;
	13'h126D: q=8'h0;
	13'h126E: q=8'hBA;
	13'h126F: q=8'h8C;
	13'h1270: q=8'hDE;
	13'h1271: q=8'hB5;
	13'h1272: q=8'h96;
	13'h1273: q=8'hC9;
	13'h1274: q=8'hA7;
	13'h1275: q=8'h0;
	13'h1276: q=8'h96;
	13'h1277: q=8'hCE;
	13'h1278: q=8'h8A;
	13'h1279: q=8'h7F;
	13'h127A: q=8'h94;
	13'h127B: q=8'hCA;
	13'h127C: q=8'hA7;
	13'h127D: q=8'h1;
	13'h127E: q=8'h96;
	13'h127F: q=8'hCB;
	13'h1280: q=8'hA7;
	13'h1281: q=8'h2;
	13'h1282: q=8'h96;
	13'h1283: q=8'hCC;
	13'h1284: q=8'hA7;
	13'h1285: q=8'h3;
	13'h1286: q=8'h96;
	13'h1287: q=8'hCD;
	13'h1288: q=8'hA7;
	13'h1289: q=8'h4;
	13'h128A: q=8'h39;
	13'h128B: q=8'h96;
	13'h128C: q=8'hDB;
	13'h128D: q=8'h97;
	13'h128E: q=8'hCE;
	13'h128F: q=8'hDE;
	13'h1290: q=8'hD6;
	13'h1291: q=8'hDF;
	13'h1292: q=8'hC9;
	13'h1293: q=8'h7F;
	13'h1294: q=8'h0;
	13'h1295: q=8'hDD;
	13'h1296: q=8'hDE;
	13'h1297: q=8'hD8;
	13'h1298: q=8'hDF;
	13'h1299: q=8'hCB;
	13'h129A: q=8'hDE;
	13'h129B: q=8'hD9;
	13'h129C: q=8'hDF;
	13'h129D: q=8'hCC;
	13'h129E: q=8'h39;
	13'h129F: q=8'hDC;
	13'h12A0: q=8'hC9;
	13'h12A1: q=8'hDD;
	13'h12A2: q=8'hD6;
	13'h12A3: q=8'hDE;
	13'h12A4: q=8'hCB;
	13'h12A5: q=8'hDF;
	13'h12A6: q=8'hD8;
	13'h12A7: q=8'hDE;
	13'h12A8: q=8'hCD;
	13'h12A9: q=8'hDF;
	13'h12AA: q=8'hDA;
	13'h12AB: q=8'h4D;
	13'h12AC: q=8'h39;
	13'h12AD: q=8'hD6;
	13'h12AE: q=8'hC9;
	13'h12AF: q=8'h27;
	13'h12B0: q=8'h8;
	13'h12B1: q=8'hD6;
	13'h12B2: q=8'hCE;
	13'h12B3: q=8'h59;
	13'h12B4: q=8'hC6;
	13'h12B5: q=8'hFF;
	13'h12B6: q=8'h25;
	13'h12B7: q=8'h1;
	13'h12B8: q=8'h50;
	13'h12B9: q=8'h39;
	13'h12BA: q=8'h8D;
	13'h12BB: q=8'hF1;
	13'h12BC: q=8'hD7;
	13'h12BD: q=8'hCA;
	13'h12BE: q=8'h7F;
	13'h12BF: q=8'h0;
	13'h12C0: q=8'hCB;
	13'h12C1: q=8'hC6;
	13'h12C2: q=8'h88;
	13'h12C3: q=8'h96;
	13'h12C4: q=8'hCA;
	13'h12C5: q=8'h80;
	13'h12C6: q=8'h80;
	13'h12C7: q=8'hD7;
	13'h12C8: q=8'hC9;
	13'h12C9: q=8'h86;
	13'h12CA: q=8'h0;
	13'h12CB: q=8'h16;
	13'h12CC: q=8'hDD;
	13'h12CD: q=8'hCC;
	13'h12CE: q=8'h97;
	13'h12CF: q=8'hDD;
	13'h12D0: q=8'h97;
	13'h12D1: q=8'hCE;
	13'h12D2: q=8'h7E;
	13'h12D3: q=8'hEF;
	13'h12D4: q=8'hD2;
	13'h12D5: q=8'h7F;
	13'h12D6: q=8'h0;
	13'h12D7: q=8'hCE;
	13'h12D8: q=8'h39;
	13'h12D9: q=8'hE6;
	13'h12DA: q=8'h0;
	13'h12DB: q=8'h27;
	13'h12DC: q=8'hD0;
	13'h12DD: q=8'hE6;
	13'h12DE: q=8'h1;
	13'h12DF: q=8'hD8;
	13'h12E0: q=8'hCE;
	13'h12E1: q=8'h2B;
	13'h12E2: q=8'hCE;
	13'h12E3: q=8'hD6;
	13'h12E4: q=8'hC9;
	13'h12E5: q=8'hE1;
	13'h12E6: q=8'h0;
	13'h12E7: q=8'h26;
	13'h12E8: q=8'h1D;
	13'h12E9: q=8'hE6;
	13'h12EA: q=8'h1;
	13'h12EB: q=8'hCA;
	13'h12EC: q=8'h7F;
	13'h12ED: q=8'hD4;
	13'h12EE: q=8'hCA;
	13'h12EF: q=8'hE1;
	13'h12F0: q=8'h1;
	13'h12F1: q=8'h26;
	13'h12F2: q=8'h13;
	13'h12F3: q=8'hD6;
	13'h12F4: q=8'hCB;
	13'h12F5: q=8'hE1;
	13'h12F6: q=8'h2;
	13'h12F7: q=8'h26;
	13'h12F8: q=8'hD;
	13'h12F9: q=8'hD6;
	13'h12FA: q=8'hCC;
	13'h12FB: q=8'hE1;
	13'h12FC: q=8'h3;
	13'h12FD: q=8'h26;
	13'h12FE: q=8'h7;
	13'h12FF: q=8'hD6;
	13'h1300: q=8'hCD;
	13'h1301: q=8'hE0;
	13'h1302: q=8'h4;
	13'h1303: q=8'h26;
	13'h1304: q=8'h1;
	13'h1305: q=8'h39;
	13'h1306: q=8'h56;
	13'h1307: q=8'hD8;
	13'h1308: q=8'hCE;
	13'h1309: q=8'h20;
	13'h130A: q=8'hA8;
	13'h130B: q=8'hD6;
	13'h130C: q=8'hC9;
	13'h130D: q=8'h27;
	13'h130E: q=8'h41;
	13'h130F: q=8'hC0;
	13'h1310: q=8'hA0;
	13'h1311: q=8'h96;
	13'h1312: q=8'hCE;
	13'h1313: q=8'h2A;
	13'h1314: q=8'h6;
	13'h1315: q=8'h73;
	13'h1316: q=8'h0;
	13'h1317: q=8'hD5;
	13'h1318: q=8'hBD;
	13'h1319: q=8'hF0;
	13'h131A: q=8'h3F;
	13'h131B: q=8'hCE;
	13'h131C: q=8'h0;
	13'h131D: q=8'hC9;
	13'h131E: q=8'hC1;
	13'h131F: q=8'hF8;
	13'h1320: q=8'h2E;
	13'h1321: q=8'h7;
	13'h1322: q=8'hBD;
	13'h1323: q=8'hF0;
	13'h1324: q=8'h74;
	13'h1325: q=8'h7F;
	13'h1326: q=8'h0;
	13'h1327: q=8'hD5;
	13'h1328: q=8'h39;
	13'h1329: q=8'h7F;
	13'h132A: q=8'h0;
	13'h132B: q=8'hD5;
	13'h132C: q=8'h96;
	13'h132D: q=8'hCE;
	13'h132E: q=8'h49;
	13'h132F: q=8'h76;
	13'h1330: q=8'h0;
	13'h1331: q=8'hCA;
	13'h1332: q=8'h7E;
	13'h1333: q=8'hF0;
	13'h1334: q=8'h80;
	13'h1335: q=8'hD6;
	13'h1336: q=8'hC9;
	13'h1337: q=8'hC1;
	13'h1338: q=8'hA0;
	13'h1339: q=8'h24;
	13'h133A: q=8'h1D;
	13'h133B: q=8'h8D;
	13'h133C: q=8'hCE;
	13'h133D: q=8'hD7;
	13'h133E: q=8'hDD;
	13'h133F: q=8'h96;
	13'h1340: q=8'hCE;
	13'h1341: q=8'hD7;
	13'h1342: q=8'hCE;
	13'h1343: q=8'h80;
	13'h1344: q=8'h80;
	13'h1345: q=8'h86;
	13'h1346: q=8'hA0;
	13'h1347: q=8'h97;
	13'h1348: q=8'hC9;
	13'h1349: q=8'h96;
	13'h134A: q=8'hCD;
	13'h134B: q=8'h97;
	13'h134C: q=8'h80;
	13'h134D: q=8'h7E;
	13'h134E: q=8'hEF;
	13'h134F: q=8'hD2;
	13'h1350: q=8'hD7;
	13'h1351: q=8'hCA;
	13'h1352: q=8'hD7;
	13'h1353: q=8'hCB;
	13'h1354: q=8'hD7;
	13'h1355: q=8'hCC;
	13'h1356: q=8'hD7;
	13'h1357: q=8'hCD;
	13'h1358: q=8'h39;
	13'h1359: q=8'hBD;
	13'h135A: q=8'h42;
	13'h135B: q=8'h9D;
	13'h135C: q=8'hCE;
	13'h135D: q=8'h0;
	13'h135E: q=8'h0;
	13'h135F: q=8'hDF;
	13'h1360: q=8'hCE;
	13'h1361: q=8'hDF;
	13'h1362: q=8'hC9;
	13'h1363: q=8'hDF;
	13'h1364: q=8'hCB;
	13'h1365: q=8'hDF;
	13'h1366: q=8'hCC;
	13'h1367: q=8'hDF;
	13'h1368: q=8'hC1;
	13'h1369: q=8'hDF;
	13'h136A: q=8'hBF;
	13'h136B: q=8'h25;
	13'h136C: q=8'h6B;
	13'h136D: q=8'h81;
	13'h136E: q=8'h2D;
	13'h136F: q=8'h26;
	13'h1370: q=8'h5;
	13'h1371: q=8'h73;
	13'h1372: q=8'h0;
	13'h1373: q=8'hCF;
	13'h1374: q=8'h20;
	13'h1375: q=8'h4;
	13'h1376: q=8'h81;
	13'h1377: q=8'h2B;
	13'h1378: q=8'h26;
	13'h1379: q=8'h5;
	13'h137A: q=8'hBD;
	13'h137B: q=8'h0;
	13'h137C: q=8'hEB;
	13'h137D: q=8'h25;
	13'h137E: q=8'h59;
	13'h137F: q=8'h81;
	13'h1380: q=8'h2E;
	13'h1381: q=8'h27;
	13'h1382: q=8'h2D;
	13'h1383: q=8'h81;
	13'h1384: q=8'h45;
	13'h1385: q=8'h26;
	13'h1386: q=8'h2E;
	13'h1387: q=8'hBD;
	13'h1388: q=8'h0;
	13'h1389: q=8'hEB;
	13'h138A: q=8'h25;
	13'h138B: q=8'h69;
	13'h138C: q=8'h81;
	13'h138D: q=8'hA8;
	13'h138E: q=8'h27;
	13'h138F: q=8'hE;
	13'h1390: q=8'h81;
	13'h1391: q=8'h2D;
	13'h1392: q=8'h27;
	13'h1393: q=8'hA;
	13'h1394: q=8'h81;
	13'h1395: q=8'hA7;
	13'h1396: q=8'h27;
	13'h1397: q=8'h9;
	13'h1398: q=8'h81;
	13'h1399: q=8'h2B;
	13'h139A: q=8'h27;
	13'h139B: q=8'h5;
	13'h139C: q=8'h20;
	13'h139D: q=8'h8;
	13'h139E: q=8'h73;
	13'h139F: q=8'h0;
	13'h13A0: q=8'hC2;
	13'h13A1: q=8'hBD;
	13'h13A2: q=8'h0;
	13'h13A3: q=8'hEB;
	13'h13A4: q=8'h25;
	13'h13A5: q=8'h4F;
	13'h13A6: q=8'h7D;
	13'h13A7: q=8'h0;
	13'h13A8: q=8'hC2;
	13'h13A9: q=8'h27;
	13'h13AA: q=8'hA;
	13'h13AB: q=8'h70;
	13'h13AC: q=8'h0;
	13'h13AD: q=8'hC1;
	13'h13AE: q=8'h20;
	13'h13AF: q=8'h5;
	13'h13B0: q=8'h73;
	13'h13B1: q=8'h0;
	13'h13B2: q=8'hC0;
	13'h13B3: q=8'h26;
	13'h13B4: q=8'hC5;
	13'h13B5: q=8'h96;
	13'h13B6: q=8'hC1;
	13'h13B7: q=8'h90;
	13'h13B8: q=8'hBF;
	13'h13B9: q=8'h97;
	13'h13BA: q=8'hC1;
	13'h13BB: q=8'h27;
	13'h13BC: q=8'h14;
	13'h13BD: q=8'h2A;
	13'h13BE: q=8'hA;
	13'h13BF: q=8'hBD;
	13'h13C0: q=8'hF1;
	13'h13C1: q=8'hB9;
	13'h13C2: q=8'h7C;
	13'h13C3: q=8'h0;
	13'h13C4: q=8'hC1;
	13'h13C5: q=8'h26;
	13'h13C6: q=8'hF8;
	13'h13C7: q=8'h20;
	13'h13C8: q=8'h8;
	13'h13C9: q=8'hBD;
	13'h13CA: q=8'hF1;
	13'h13CB: q=8'h9F;
	13'h13CC: q=8'h7A;
	13'h13CD: q=8'h0;
	13'h13CE: q=8'hC1;
	13'h13CF: q=8'h26;
	13'h13D0: q=8'hF8;
	13'h13D1: q=8'h96;
	13'h13D2: q=8'hCF;
	13'h13D3: q=8'h2A;
	13'h13D4: q=8'h83;
	13'h13D5: q=8'h7E;
	13'h13D6: q=8'hF5;
	13'h13D7: q=8'h93;
	13'h13D8: q=8'hD6;
	13'h13D9: q=8'hBF;
	13'h13DA: q=8'hD0;
	13'h13DB: q=8'hC0;
	13'h13DC: q=8'hD7;
	13'h13DD: q=8'hBF;
	13'h13DE: q=8'h36;
	13'h13DF: q=8'hBD;
	13'h13E0: q=8'hF1;
	13'h13E1: q=8'h9F;
	13'h13E2: q=8'h33;
	13'h13E3: q=8'hC0;
	13'h13E4: q=8'h30;
	13'h13E5: q=8'h8D;
	13'h13E6: q=8'h2;
	13'h13E7: q=8'h20;
	13'h13E8: q=8'h91;
	13'h13E9: q=8'hBD;
	13'h13EA: q=8'hF2;
	13'h13EB: q=8'h6C;
	13'h13EC: q=8'hBD;
	13'h13ED: q=8'hF2;
	13'h13EE: q=8'hBC;
	13'h13EF: q=8'hCE;
	13'h13F0: q=8'h0;
	13'h13F1: q=8'hBA;
	13'h13F2: q=8'h7E;
	13'h13F3: q=8'hEF;
	13'h13F4: q=8'h7D;
	13'h13F5: q=8'hD6;
	13'h13F6: q=8'hC1;
	13'h13F7: q=8'h58;
	13'h13F8: q=8'h58;
	13'h13F9: q=8'hDB;
	13'h13FA: q=8'hC1;
	13'h13FB: q=8'h58;
	13'h13FC: q=8'h80;
	13'h13FD: q=8'h30;
	13'h13FE: q=8'h1B;
	13'h13FF: q=8'h97;
	13'h1400: q=8'hC1;
	13'h1401: q=8'h20;
	13'h1402: q=8'h9E;
	13'h1403: q=8'h9B;
	13'h1404: q=8'h3E;
	13'h1405: q=8'hBC;
	13'h1406: q=8'h1F;
	13'h1407: q=8'hFD;
	13'h1408: q=8'h9E;
	13'h1409: q=8'h6E;
	13'h140A: q=8'h6B;
	13'h140B: q=8'h27;
	13'h140C: q=8'hFD;
	13'h140D: q=8'h9E;
	13'h140E: q=8'h6E;
	13'h140F: q=8'h6B;
	13'h1410: q=8'h28;
	13'h1411: q=8'h0;
	13'h1412: q=8'hCE;
	13'h1413: q=8'hE1;
	13'h1414: q=8'hB6;
	13'h1415: q=8'h8D;
	13'h1416: q=8'hC;
	13'h1417: q=8'hDC;
	13'h1418: q=8'hE2;
	13'h1419: q=8'hDD;
	13'h141A: q=8'hCA;
	13'h141B: q=8'hC6;
	13'h141C: q=8'h90;
	13'h141D: q=8'hD;
	13'h141E: q=8'hBD;
	13'h141F: q=8'hF2;
	13'h1420: q=8'hC7;
	13'h1421: q=8'h8D;
	13'h1422: q=8'h3;
	13'h1423: q=8'h7E;
	13'h1424: q=8'hE7;
	13'h1425: q=8'hA8;
	13'h1426: q=8'hCE;
	13'h1427: q=8'h43;
	13'h1428: q=8'h35;
	13'h1429: q=8'h86;
	13'h142A: q=8'h20;
	13'h142B: q=8'hD6;
	13'h142C: q=8'hCE;
	13'h142D: q=8'h2A;
	13'h142E: q=8'h2;
	13'h142F: q=8'h86;
	13'h1430: q=8'h2D;
	13'h1431: q=8'hA7;
	13'h1432: q=8'h0;
	13'h1433: q=8'h97;
	13'h1434: q=8'hCE;
	13'h1435: q=8'hDF;
	13'h1436: q=8'hDE;
	13'h1437: q=8'h8;
	13'h1438: q=8'h86;
	13'h1439: q=8'h30;
	13'h143A: q=8'hD6;
	13'h143B: q=8'hC9;
	13'h143C: q=8'h26;
	13'h143D: q=8'h3;
	13'h143E: q=8'h7E;
	13'h143F: q=8'hF5;
	13'h1440: q=8'h1C;
	13'h1441: q=8'h4F;
	13'h1442: q=8'hC1;
	13'h1443: q=8'h80;
	13'h1444: q=8'h22;
	13'h1445: q=8'h8;
	13'h1446: q=8'hCE;
	13'h1447: q=8'hF4;
	13'h1448: q=8'hD;
	13'h1449: q=8'hBD;
	13'h144A: q=8'hF0;
	13'h144B: q=8'hEF;
	13'h144C: q=8'h86;
	13'h144D: q=8'hF7;
	13'h144E: q=8'h97;
	13'h144F: q=8'hBF;
	13'h1450: q=8'hCE;
	13'h1451: q=8'hF4;
	13'h1452: q=8'h8;
	13'h1453: q=8'hBD;
	13'h1454: q=8'hF2;
	13'h1455: q=8'hE3;
	13'h1456: q=8'h2E;
	13'h1457: q=8'h10;
	13'h1458: q=8'hCE;
	13'h1459: q=8'hF4;
	13'h145A: q=8'h3;
	13'h145B: q=8'hBD;
	13'h145C: q=8'hF2;
	13'h145D: q=8'hE3;
	13'h145E: q=8'h2E;
	13'h145F: q=8'h10;
	13'h1460: q=8'hBD;
	13'h1461: q=8'hF1;
	13'h1462: q=8'h9F;
	13'h1463: q=8'h7A;
	13'h1464: q=8'h0;
	13'h1465: q=8'hBF;
	13'h1466: q=8'h20;
	13'h1467: q=8'hF0;
	13'h1468: q=8'hBD;
	13'h1469: q=8'hF1;
	13'h146A: q=8'hB9;
	13'h146B: q=8'h7C;
	13'h146C: q=8'h0;
	13'h146D: q=8'hBF;
	13'h146E: q=8'h20;
	13'h146F: q=8'hE0;
	13'h1470: q=8'hBD;
	13'h1471: q=8'hEF;
	13'h1472: q=8'h6D;
	13'h1473: q=8'hBD;
	13'h1474: q=8'hF3;
	13'h1475: q=8'hB;
	13'h1476: q=8'hC6;
	13'h1477: q=8'h1;
	13'h1478: q=8'h96;
	13'h1479: q=8'hBF;
	13'h147A: q=8'h8B;
	13'h147B: q=8'hA;
	13'h147C: q=8'h2B;
	13'h147D: q=8'h8;
	13'h147E: q=8'h81;
	13'h147F: q=8'hB;
	13'h1480: q=8'h24;
	13'h1481: q=8'h4;
	13'h1482: q=8'h4A;
	13'h1483: q=8'h16;
	13'h1484: q=8'h86;
	13'h1485: q=8'h2;
	13'h1486: q=8'h4A;
	13'h1487: q=8'h4A;
	13'h1488: q=8'h97;
	13'h1489: q=8'hC1;
	13'h148A: q=8'hD7;
	13'h148B: q=8'hBF;
	13'h148C: q=8'h2E;
	13'h148D: q=8'h11;
	13'h148E: q=8'hDE;
	13'h148F: q=8'hDE;
	13'h1490: q=8'h86;
	13'h1491: q=8'h2E;
	13'h1492: q=8'h8;
	13'h1493: q=8'hA7;
	13'h1494: q=8'h0;
	13'h1495: q=8'h5D;
	13'h1496: q=8'h27;
	13'h1497: q=8'h5;
	13'h1498: q=8'h86;
	13'h1499: q=8'h30;
	13'h149A: q=8'h8;
	13'h149B: q=8'hA7;
	13'h149C: q=8'h0;
	13'h149D: q=8'hDF;
	13'h149E: q=8'hDE;
	13'h149F: q=8'hCE;
	13'h14A0: q=8'hF5;
	13'h14A1: q=8'h29;
	13'h14A2: q=8'hC6;
	13'h14A3: q=8'h80;
	13'h14A4: q=8'h96;
	13'h14A5: q=8'hCD;
	13'h14A6: q=8'hAB;
	13'h14A7: q=8'h3;
	13'h14A8: q=8'h97;
	13'h14A9: q=8'hCD;
	13'h14AA: q=8'h96;
	13'h14AB: q=8'hCC;
	13'h14AC: q=8'hA9;
	13'h14AD: q=8'h2;
	13'h14AE: q=8'h97;
	13'h14AF: q=8'hCC;
	13'h14B0: q=8'h96;
	13'h14B1: q=8'hCB;
	13'h14B2: q=8'hA9;
	13'h14B3: q=8'h1;
	13'h14B4: q=8'h97;
	13'h14B5: q=8'hCB;
	13'h14B6: q=8'h96;
	13'h14B7: q=8'hCA;
	13'h14B8: q=8'hA9;
	13'h14B9: q=8'h0;
	13'h14BA: q=8'h97;
	13'h14BB: q=8'hCA;
	13'h14BC: q=8'h5C;
	13'h14BD: q=8'h56;
	13'h14BE: q=8'h59;
	13'h14BF: q=8'h28;
	13'h14C0: q=8'hE3;
	13'h14C1: q=8'h24;
	13'h14C2: q=8'h3;
	13'h14C3: q=8'hC0;
	13'h14C4: q=8'hB;
	13'h14C5: q=8'h50;
	13'h14C6: q=8'hCB;
	13'h14C7: q=8'h2F;
	13'h14C8: q=8'h8;
	13'h14C9: q=8'h8;
	13'h14CA: q=8'h8;
	13'h14CB: q=8'h8;
	13'h14CC: q=8'hDF;
	13'h14CD: q=8'hB3;
	13'h14CE: q=8'hDE;
	13'h14CF: q=8'hDE;
	13'h14D0: q=8'h8;
	13'h14D1: q=8'h17;
	13'h14D2: q=8'h84;
	13'h14D3: q=8'h7F;
	13'h14D4: q=8'hA7;
	13'h14D5: q=8'h0;
	13'h14D6: q=8'h7A;
	13'h14D7: q=8'h0;
	13'h14D8: q=8'hBF;
	13'h14D9: q=8'h26;
	13'h14DA: q=8'h5;
	13'h14DB: q=8'h86;
	13'h14DC: q=8'h2E;
	13'h14DD: q=8'h8;
	13'h14DE: q=8'hA7;
	13'h14DF: q=8'h0;
	13'h14E0: q=8'hDF;
	13'h14E1: q=8'hDE;
	13'h14E2: q=8'hDE;
	13'h14E3: q=8'hB3;
	13'h14E4: q=8'h53;
	13'h14E5: q=8'hC4;
	13'h14E6: q=8'h80;
	13'h14E7: q=8'h8C;
	13'h14E8: q=8'hF5;
	13'h14E9: q=8'h4D;
	13'h14EA: q=8'h26;
	13'h14EB: q=8'hB8;
	13'h14EC: q=8'hDE;
	13'h14ED: q=8'hDE;
	13'h14EE: q=8'hA6;
	13'h14EF: q=8'h0;
	13'h14F0: q=8'h9;
	13'h14F1: q=8'h81;
	13'h14F2: q=8'h30;
	13'h14F3: q=8'h27;
	13'h14F4: q=8'hF9;
	13'h14F5: q=8'h81;
	13'h14F6: q=8'h2E;
	13'h14F7: q=8'h27;
	13'h14F8: q=8'h1;
	13'h14F9: q=8'h8;
	13'h14FA: q=8'h86;
	13'h14FB: q=8'h2B;
	13'h14FC: q=8'hD6;
	13'h14FD: q=8'hC1;
	13'h14FE: q=8'h27;
	13'h14FF: q=8'h1E;
	13'h1500: q=8'h2A;
	13'h1501: q=8'h3;
	13'h1502: q=8'h86;
	13'h1503: q=8'h2D;
	13'h1504: q=8'h50;
	13'h1505: q=8'hA7;
	13'h1506: q=8'h2;
	13'h1507: q=8'h86;
	13'h1508: q=8'h45;
	13'h1509: q=8'hA7;
	13'h150A: q=8'h1;
	13'h150B: q=8'h86;
	13'h150C: q=8'h2F;
	13'h150D: q=8'h4C;
	13'h150E: q=8'hC0;
	13'h150F: q=8'hA;
	13'h1510: q=8'h24;
	13'h1511: q=8'hFB;
	13'h1512: q=8'hCB;
	13'h1513: q=8'h3A;
	13'h1514: q=8'hA7;
	13'h1515: q=8'h3;
	13'h1516: q=8'hE7;
	13'h1517: q=8'h4;
	13'h1518: q=8'h6F;
	13'h1519: q=8'h5;
	13'h151A: q=8'h20;
	13'h151B: q=8'h4;
	13'h151C: q=8'hA7;
	13'h151D: q=8'h0;
	13'h151E: q=8'h6F;
	13'h151F: q=8'h1;
	13'h1520: q=8'hCE;
	13'h1521: q=8'h43;
	13'h1522: q=8'h35;
	13'h1523: q=8'h39;
	13'h1524: q=8'h80;
	13'h1525: q=8'h0;
	13'h1526: q=8'h0;
	13'h1527: q=8'h0;
	13'h1528: q=8'h0;
	13'h1529: q=8'hFA;
	13'h152A: q=8'hA;
	13'h152B: q=8'h1F;
	13'h152C: q=8'h0;
	13'h152D: q=8'h0;
	13'h152E: q=8'h98;
	13'h152F: q=8'h96;
	13'h1530: q=8'h80;
	13'h1531: q=8'hFF;
	13'h1532: q=8'hF0;
	13'h1533: q=8'hBD;
	13'h1534: q=8'hC0;
	13'h1535: q=8'h0;
	13'h1536: q=8'h1;
	13'h1537: q=8'h86;
	13'h1538: q=8'hA0;
	13'h1539: q=8'hFF;
	13'h153A: q=8'hFF;
	13'h153B: q=8'hD8;
	13'h153C: q=8'hF0;
	13'h153D: q=8'h0;
	13'h153E: q=8'h0;
	13'h153F: q=8'h3;
	13'h1540: q=8'hE8;
	13'h1541: q=8'hFF;
	13'h1542: q=8'hFF;
	13'h1543: q=8'hFF;
	13'h1544: q=8'h9C;
	13'h1545: q=8'h0;
	13'h1546: q=8'h0;
	13'h1547: q=8'h0;
	13'h1548: q=8'hA;
	13'h1549: q=8'hFF;
	13'h154A: q=8'hFF;
	13'h154B: q=8'hFF;
	13'h154C: q=8'hFF;
	13'h154D: q=8'hBD;
	13'h154E: q=8'hF2;
	13'h154F: q=8'h9F;
	13'h1550: q=8'hCE;
	13'h1551: q=8'hF5;
	13'h1552: q=8'h24;
	13'h1553: q=8'hBD;
	13'h1554: q=8'hF2;
	13'h1555: q=8'h51;
	13'h1556: q=8'h27;
	13'h1557: q=8'h71;
	13'h1558: q=8'h4D;
	13'h1559: q=8'h26;
	13'h155A: q=8'hA;
	13'h155B: q=8'h96;
	13'h155C: q=8'hCE;
	13'h155D: q=8'h2A;
	13'h155E: q=8'h3;
	13'h155F: q=8'h7E;
	13'h1560: q=8'hF2;
	13'h1561: q=8'h43;
	13'h1562: q=8'h7E;
	13'h1563: q=8'hEF;
	13'h1564: q=8'hF5;
	13'h1565: q=8'hCE;
	13'h1566: q=8'h0;
	13'h1567: q=8'hC4;
	13'h1568: q=8'hBD;
	13'h1569: q=8'hF2;
	13'h156A: q=8'h72;
	13'h156B: q=8'h5F;
	13'h156C: q=8'h96;
	13'h156D: q=8'hDB;
	13'h156E: q=8'h2A;
	13'h156F: q=8'h10;
	13'h1570: q=8'hBD;
	13'h1571: q=8'hF3;
	13'h1572: q=8'h35;
	13'h1573: q=8'hCE;
	13'h1574: q=8'h0;
	13'h1575: q=8'hC4;
	13'h1576: q=8'h96;
	13'h1577: q=8'hDB;
	13'h1578: q=8'hBD;
	13'h1579: q=8'hF2;
	13'h157A: q=8'hE3;
	13'h157B: q=8'h26;
	13'h157C: q=8'h3;
	13'h157D: q=8'h43;
	13'h157E: q=8'hD6;
	13'h157F: q=8'h80;
	13'h1580: q=8'hBD;
	13'h1581: q=8'hF2;
	13'h1582: q=8'h8D;
	13'h1583: q=8'h37;
	13'h1584: q=8'hBD;
	13'h1585: q=8'hF0;
	13'h1586: q=8'hB9;
	13'h1587: q=8'hCE;
	13'h1588: q=8'h0;
	13'h1589: q=8'hC4;
	13'h158A: q=8'hBD;
	13'h158B: q=8'hF0;
	13'h158C: q=8'hEF;
	13'h158D: q=8'h8D;
	13'h158E: q=8'h3A;
	13'h158F: q=8'h32;
	13'h1590: q=8'h46;
	13'h1591: q=8'h24;
	13'h1592: q=8'h90;
	13'h1593: q=8'h96;
	13'h1594: q=8'hC9;
	13'h1595: q=8'h27;
	13'h1596: q=8'h3;
	13'h1597: q=8'h73;
	13'h1598: q=8'h0;
	13'h1599: q=8'hCE;
	13'h159A: q=8'h39;
	13'h159B: q=8'h81;
	13'h159C: q=8'h38;
	13'h159D: q=8'hAA;
	13'h159E: q=8'h3B;
	13'h159F: q=8'h29;
	13'h15A0: q=8'h7;
	13'h15A1: q=8'h71;
	13'h15A2: q=8'h34;
	13'h15A3: q=8'h58;
	13'h15A4: q=8'h3E;
	13'h15A5: q=8'h56;
	13'h15A6: q=8'h74;
	13'h15A7: q=8'h16;
	13'h15A8: q=8'h7E;
	13'h15A9: q=8'hB3;
	13'h15AA: q=8'h1B;
	13'h15AB: q=8'h77;
	13'h15AC: q=8'h2F;
	13'h15AD: q=8'hEE;
	13'h15AE: q=8'hE3;
	13'h15AF: q=8'h85;
	13'h15B0: q=8'h7A;
	13'h15B1: q=8'h1D;
	13'h15B2: q=8'h84;
	13'h15B3: q=8'h1C;
	13'h15B4: q=8'h2A;
	13'h15B5: q=8'h7C;
	13'h15B6: q=8'h63;
	13'h15B7: q=8'h59;
	13'h15B8: q=8'h58;
	13'h15B9: q=8'hA;
	13'h15BA: q=8'h7E;
	13'h15BB: q=8'h75;
	13'h15BC: q=8'hFD;
	13'h15BD: q=8'hE7;
	13'h15BE: q=8'hC6;
	13'h15BF: q=8'h80;
	13'h15C0: q=8'h31;
	13'h15C1: q=8'h72;
	13'h15C2: q=8'h18;
	13'h15C3: q=8'h10;
	13'h15C4: q=8'h81;
	13'h15C5: q=8'h0;
	13'h15C6: q=8'h0;
	13'h15C7: q=8'h0;
	13'h15C8: q=8'h0;
	13'h15C9: q=8'hCE;
	13'h15CA: q=8'hF5;
	13'h15CB: q=8'h9B;
	13'h15CC: q=8'h8D;
	13'h15CD: q=8'h36;
	13'h15CE: q=8'hBD;
	13'h15CF: q=8'hF2;
	13'h15D0: q=8'h6C;
	13'h15D1: q=8'h96;
	13'h15D2: q=8'hC9;
	13'h15D3: q=8'h81;
	13'h15D4: q=8'h88;
	13'h15D5: q=8'h25;
	13'h15D6: q=8'h3;
	13'h15D7: q=8'h7E;
	13'h15D8: q=8'hF1;
	13'h15D9: q=8'h90;
	13'h15DA: q=8'hBD;
	13'h15DB: q=8'hF3;
	13'h15DC: q=8'h35;
	13'h15DD: q=8'h96;
	13'h15DE: q=8'h80;
	13'h15DF: q=8'h8B;
	13'h15E0: q=8'h81;
	13'h15E1: q=8'h27;
	13'h15E2: q=8'hF4;
	13'h15E3: q=8'h4A;
	13'h15E4: q=8'h36;
	13'h15E5: q=8'hCE;
	13'h15E6: q=8'h0;
	13'h15E7: q=8'hBA;
	13'h15E8: q=8'hBD;
	13'h15E9: q=8'hEF;
	13'h15EA: q=8'h72;
	13'h15EB: q=8'hCE;
	13'h15EC: q=8'hF5;
	13'h15ED: q=8'hA0;
	13'h15EE: q=8'h8D;
	13'h15EF: q=8'h17;
	13'h15F0: q=8'h7F;
	13'h15F1: q=8'h0;
	13'h15F2: q=8'hDC;
	13'h15F3: q=8'h32;
	13'h15F4: q=8'hBD;
	13'h15F5: q=8'hF1;
	13'h15F6: q=8'h79;
	13'h15F7: q=8'h39;
	13'h15F8: q=8'hDF;
	13'h15F9: q=8'hDE;
	13'h15FA: q=8'hBD;
	13'h15FB: q=8'hF2;
	13'h15FC: q=8'h6C;
	13'h15FD: q=8'h8D;
	13'h15FE: q=8'h5;
	13'h15FF: q=8'h8D;
	13'h1600: q=8'h8;
	13'h1601: q=8'hCE;
	13'h1602: q=8'h0;
	13'h1603: q=8'hBA;
	13'h1604: q=8'h7E;
	13'h1605: q=8'hF0;
	13'h1606: q=8'hEF;
	13'h1607: q=8'hDF;
	13'h1608: q=8'hDE;
	13'h1609: q=8'hBD;
	13'h160A: q=8'hF2;
	13'h160B: q=8'h67;
	13'h160C: q=8'hDE;
	13'h160D: q=8'hDE;
	13'h160E: q=8'hE6;
	13'h160F: q=8'h0;
	13'h1610: q=8'hD7;
	13'h1611: q=8'hCF;
	13'h1612: q=8'h8;
	13'h1613: q=8'hDF;
	13'h1614: q=8'hDE;
	13'h1615: q=8'h8D;
	13'h1616: q=8'hED;
	13'h1617: q=8'hDE;
	13'h1618: q=8'hDE;
	13'h1619: q=8'hC6;
	13'h161A: q=8'h5;
	13'h161B: q=8'h3A;
	13'h161C: q=8'hDF;
	13'h161D: q=8'hDE;
	13'h161E: q=8'hBD;
	13'h161F: q=8'hEF;
	13'h1620: q=8'h7D;
	13'h1621: q=8'hCE;
	13'h1622: q=8'h0;
	13'h1623: q=8'hBF;
	13'h1624: q=8'h7A;
	13'h1625: q=8'h0;
	13'h1626: q=8'hCF;
	13'h1627: q=8'h26;
	13'h1628: q=8'hEC;
	13'h1629: q=8'h39;
	13'h162A: q=8'hBD;
	13'h162B: q=8'hF2;
	13'h162C: q=8'hAD;
	13'h162D: q=8'h2B;
	13'h162E: q=8'h21;
	13'h162F: q=8'h27;
	13'h1630: q=8'h15;
	13'h1631: q=8'h8D;
	13'h1632: q=8'h10;
	13'h1633: q=8'hBD;
	13'h1634: q=8'hF2;
	13'h1635: q=8'h6C;
	13'h1636: q=8'h8D;
	13'h1637: q=8'hE;
	13'h1638: q=8'hCE;
	13'h1639: q=8'h0;
	13'h163A: q=8'hBA;
	13'h163B: q=8'h8D;
	13'h163C: q=8'hC7;
	13'h163D: q=8'hCE;
	13'h163E: q=8'hF0;
	13'h163F: q=8'h8B;
	13'h1640: q=8'hBD;
	13'h1641: q=8'hEF;
	13'h1642: q=8'h7D;
	13'h1643: q=8'h7E;
	13'h1644: q=8'hF3;
	13'h1645: q=8'h35;
	13'h1646: q=8'hFE;
	13'h1647: q=8'h42;
	13'h1648: q=8'h18;
	13'h1649: q=8'hDF;
	13'h164A: q=8'hCA;
	13'h164B: q=8'hFE;
	13'h164C: q=8'h42;
	13'h164D: q=8'h1A;
	13'h164E: q=8'hDF;
	13'h164F: q=8'hCC;
	13'h1650: q=8'hFE;
	13'h1651: q=8'hF6;
	13'h1652: q=8'h82;
	13'h1653: q=8'hDF;
	13'h1654: q=8'hD7;
	13'h1655: q=8'hFE;
	13'h1656: q=8'hF6;
	13'h1657: q=8'h84;
	13'h1658: q=8'hDF;
	13'h1659: q=8'hD9;
	13'h165A: q=8'hBD;
	13'h165B: q=8'hF0;
	13'h165C: q=8'hF6;
	13'h165D: q=8'hFC;
	13'h165E: q=8'h42;
	13'h165F: q=8'h54;
	13'h1660: q=8'hC3;
	13'h1661: q=8'h65;
	13'h1662: q=8'h8B;
	13'h1663: q=8'hFD;
	13'h1664: q=8'h42;
	13'h1665: q=8'h1A;
	13'h1666: q=8'hDD;
	13'h1667: q=8'hCC;
	13'h1668: q=8'hFC;
	13'h1669: q=8'h42;
	13'h166A: q=8'h52;
	13'h166B: q=8'hC9;
	13'h166C: q=8'hB0;
	13'h166D: q=8'h89;
	13'h166E: q=8'h5;
	13'h166F: q=8'hFD;
	13'h1670: q=8'h42;
	13'h1671: q=8'h18;
	13'h1672: q=8'hDD;
	13'h1673: q=8'hCA;
	13'h1674: q=8'h7F;
	13'h1675: q=8'h0;
	13'h1676: q=8'hCE;
	13'h1677: q=8'h86;
	13'h1678: q=8'h80;
	13'h1679: q=8'h97;
	13'h167A: q=8'hC9;
	13'h167B: q=8'h96;
	13'h167C: q=8'h8F;
	13'h167D: q=8'h97;
	13'h167E: q=8'hDD;
	13'h167F: q=8'h7E;
	13'h1680: q=8'hEF;
	13'h1681: q=8'hD6;
	13'h1682: q=8'h40;
	13'h1683: q=8'hE6;
	13'h1684: q=8'h4D;
	13'h1685: q=8'hAB;
	13'h1686: q=8'hCE;
	13'h1687: q=8'hF6;
	13'h1688: q=8'hF6;
	13'h1689: q=8'hBD;
	13'h168A: q=8'hEF;
	13'h168B: q=8'h7D;
	13'h168C: q=8'hBD;
	13'h168D: q=8'hF2;
	13'h168E: q=8'h9F;
	13'h168F: q=8'hCE;
	13'h1690: q=8'hF6;
	13'h1691: q=8'hFB;
	13'h1692: q=8'hD6;
	13'h1693: q=8'hDB;
	13'h1694: q=8'hBD;
	13'h1695: q=8'hF1;
	13'h1696: q=8'hC0;
	13'h1697: q=8'hBD;
	13'h1698: q=8'hF2;
	13'h1699: q=8'h9F;
	13'h169A: q=8'hBD;
	13'h169B: q=8'hF3;
	13'h169C: q=8'h35;
	13'h169D: q=8'h7F;
	13'h169E: q=8'h0;
	13'h169F: q=8'hDC;
	13'h16A0: q=8'h96;
	13'h16A1: q=8'hD6;
	13'h16A2: q=8'hD6;
	13'h16A3: q=8'hC9;
	13'h16A4: q=8'hBD;
	13'h16A5: q=8'hEF;
	13'h16A6: q=8'h75;
	13'h16A7: q=8'hCE;
	13'h16A8: q=8'hF7;
	13'h16A9: q=8'h0;
	13'h16AA: q=8'hBD;
	13'h16AB: q=8'hEF;
	13'h16AC: q=8'h72;
	13'h16AD: q=8'h96;
	13'h16AE: q=8'hCE;
	13'h16AF: q=8'h36;
	13'h16B0: q=8'h2A;
	13'h16B1: q=8'hA;
	13'h16B2: q=8'hBD;
	13'h16B3: q=8'hEF;
	13'h16B4: q=8'h6D;
	13'h16B5: q=8'h96;
	13'h16B6: q=8'hCE;
	13'h16B7: q=8'h2B;
	13'h16B8: q=8'h6;
	13'h16B9: q=8'h73;
	13'h16BA: q=8'h0;
	13'h16BB: q=8'h88;
	13'h16BC: q=8'hBD;
	13'h16BD: q=8'hF5;
	13'h16BE: q=8'h93;
	13'h16BF: q=8'hCE;
	13'h16C0: q=8'hF7;
	13'h16C1: q=8'h0;
	13'h16C2: q=8'hBD;
	13'h16C3: q=8'hEF;
	13'h16C4: q=8'h7D;
	13'h16C5: q=8'h32;
	13'h16C6: q=8'h4D;
	13'h16C7: q=8'h2A;
	13'h16C8: q=8'h3;
	13'h16C9: q=8'hBD;
	13'h16CA: q=8'hF5;
	13'h16CB: q=8'h93;
	13'h16CC: q=8'hCE;
	13'h16CD: q=8'hF7;
	13'h16CE: q=8'h5;
	13'h16CF: q=8'h7E;
	13'h16D0: q=8'hF5;
	13'h16D1: q=8'hF8;
	13'h16D2: q=8'hBD;
	13'h16D3: q=8'hF2;
	13'h16D4: q=8'h6C;
	13'h16D5: q=8'h7F;
	13'h16D6: q=8'h0;
	13'h16D7: q=8'h88;
	13'h16D8: q=8'h8D;
	13'h16D9: q=8'hB2;
	13'h16DA: q=8'hCE;
	13'h16DB: q=8'h0;
	13'h16DC: q=8'hC4;
	13'h16DD: q=8'hBD;
	13'h16DE: q=8'hF2;
	13'h16DF: q=8'h72;
	13'h16E0: q=8'hCE;
	13'h16E1: q=8'h0;
	13'h16E2: q=8'hBA;
	13'h16E3: q=8'hBD;
	13'h16E4: q=8'hF2;
	13'h16E5: q=8'h51;
	13'h16E6: q=8'h7F;
	13'h16E7: q=8'h0;
	13'h16E8: q=8'hCE;
	13'h16E9: q=8'h96;
	13'h16EA: q=8'h88;
	13'h16EB: q=8'h8D;
	13'h16EC: q=8'h6;
	13'h16ED: q=8'hCE;
	13'h16EE: q=8'h0;
	13'h16EF: q=8'hC4;
	13'h16F0: q=8'h7E;
	13'h16F1: q=8'hF1;
	13'h16F2: q=8'hC6;
	13'h16F3: q=8'h36;
	13'h16F4: q=8'h20;
	13'h16F5: q=8'hC6;
	13'h16F6: q=8'h81;
	13'h16F7: q=8'h49;
	13'h16F8: q=8'hF;
	13'h16F9: q=8'hDA;
	13'h16FA: q=8'hA2;
	13'h16FB: q=8'h83;
	13'h16FC: q=8'h49;
	13'h16FD: q=8'hF;
	13'h16FE: q=8'hDA;
	13'h16FF: q=8'hA2;
	13'h1700: q=8'h7F;
	13'h1701: q=8'h0;
	13'h1702: q=8'h0;
	13'h1703: q=8'h0;
	13'h1704: q=8'h0;
	13'h1705: q=8'h5;
	13'h1706: q=8'h84;
	13'h1707: q=8'hE6;
	13'h1708: q=8'h1A;
	13'h1709: q=8'h2D;
	13'h170A: q=8'h1B;
	13'h170B: q=8'h86;
	13'h170C: q=8'h28;
	13'h170D: q=8'h7;
	13'h170E: q=8'hFB;
	13'h170F: q=8'hF8;
	13'h1710: q=8'h87;
	13'h1711: q=8'h99;
	13'h1712: q=8'h68;
	13'h1713: q=8'h89;
	13'h1714: q=8'h1;
	13'h1715: q=8'h87;
	13'h1716: q=8'h23;
	13'h1717: q=8'h35;
	13'h1718: q=8'hDF;
	13'h1719: q=8'hE1;
	13'h171A: q=8'h86;
	13'h171B: q=8'hA5;
	13'h171C: q=8'h5D;
	13'h171D: q=8'hE7;
	13'h171E: q=8'h28;
	13'h171F: q=8'h83;
	13'h1720: q=8'h49;
	13'h1721: q=8'hF;
	13'h1722: q=8'hDA;
	13'h1723: q=8'hA2;
	13'h1724: q=8'hA1;
	13'h1725: q=8'h54;
	13'h1726: q=8'h46;
	13'h1727: q=8'h8F;
	13'h1728: q=8'h13;
	13'h1729: q=8'h8F;
	13'h172A: q=8'h52;
	13'h172B: q=8'h43;
	13'h172C: q=8'h89;
	13'h172D: q=8'hCD;
	13'h172E: q=8'h86;
	13'h172F: q=8'hFF;
	13'h1730: q=8'h97;
	13'h1731: q=8'h0;
	13'h1732: q=8'h86;
	13'h1733: q=8'h1;
	13'h1734: q=8'h97;
	13'h1735: q=8'h1;
	13'h1736: q=8'h86;
	13'h1737: q=8'h1;
	13'h1738: q=8'h97;
	13'h1739: q=8'h3;
	13'h173A: q=8'h96;
	13'h173B: q=8'hEA;
	13'h173C: q=8'h81;
	13'h173D: q=8'h55;
	13'h173E: q=8'h26;
	13'h173F: q=8'hA;
	13'h1740: q=8'hFE;
	13'h1741: q=8'h42;
	13'h1742: q=8'h21;
	13'h1743: q=8'hA6;
	13'h1744: q=8'h0;
	13'h1745: q=8'h4A;
	13'h1746: q=8'h26;
	13'h1747: q=8'h2;
	13'h1748: q=8'h6E;
	13'h1749: q=8'h0;
	13'h174A: q=8'hCE;
	13'h174B: q=8'h0;
	13'h174C: q=8'h80;
	13'h174D: q=8'h6F;
	13'h174E: q=8'h0;
	13'h174F: q=8'h8;
	13'h1750: q=8'h8C;
	13'h1751: q=8'h1;
	13'h1752: q=8'h0;
	13'h1753: q=8'h26;
	13'h1754: q=8'hF8;
	13'h1755: q=8'hCE;
	13'h1756: q=8'h41;
	13'h1757: q=8'hFD;
	13'h1758: q=8'h8;
	13'h1759: q=8'hA6;
	13'h175A: q=8'h2;
	13'h175B: q=8'h63;
	13'h175C: q=8'h2;
	13'h175D: q=8'hE6;
	13'h175E: q=8'h2;
	13'h175F: q=8'h6F;
	13'h1760: q=8'h2;
	13'h1761: q=8'h43;
	13'h1762: q=8'h11;
	13'h1763: q=8'h27;
	13'h1764: q=8'hF3;
	13'h1765: q=8'hFF;
	13'h1766: q=8'h42;
	13'h1767: q=8'h50;
	13'h1768: q=8'hDF;
	13'h1769: q=8'hA1;
	13'h176A: q=8'hDF;
	13'h176B: q=8'h9D;
	13'h176C: q=8'hDC;
	13'h176D: q=8'h9D;
	13'h176E: q=8'h83;
	13'h176F: q=8'h0;
	13'h1770: q=8'h64;
	13'h1771: q=8'hDD;
	13'h1772: q=8'h9B;
	13'h1773: q=8'h9E;
	13'h1774: q=8'h9B;
	13'h1775: q=8'hCE;
	13'h1776: q=8'hF7;
	13'h1777: q=8'hCF;
	13'h1778: q=8'hCC;
	13'h1779: q=8'h0;
	13'h177A: q=8'hEB;
	13'h177B: q=8'h8D;
	13'h177C: q=8'h30;
	13'h177D: q=8'hCE;
	13'h177E: q=8'hF7;
	13'h177F: q=8'hDE;
	13'h1780: q=8'hCC;
	13'h1781: q=8'h42;
	13'h1782: q=8'h0;
	13'h1783: q=8'h8D;
	13'h1784: q=8'h28;
	13'h1785: q=8'h86;
	13'h1786: q=8'h39;
	13'h1787: q=8'hCE;
	13'h1788: q=8'h42;
	13'h1789: q=8'h85;
	13'h178A: q=8'hA7;
	13'h178B: q=8'h0;
	13'h178C: q=8'h8;
	13'h178D: q=8'h8C;
	13'h178E: q=8'h42;
	13'h178F: q=8'hAF;
	13'h1790: q=8'h26;
	13'h1791: q=8'hF8;
	13'h1792: q=8'h73;
	13'h1793: q=8'h42;
	13'h1794: q=8'hAF;
	13'h1795: q=8'hCE;
	13'h1796: q=8'h43;
	13'h1797: q=8'h46;
	13'h1798: q=8'hDF;
	13'h1799: q=8'h93;
	13'h179A: q=8'hBD;
	13'h179B: q=8'hE3;
	13'h179C: q=8'hCF;
	13'h179D: q=8'hBD;
	13'h179E: q=8'hFB;
	13'h179F: q=8'hD4;
	13'h17A0: q=8'hCE;
	13'h17A1: q=8'hF8;
	13'h17A2: q=8'hF;
	13'h17A3: q=8'hBD;
	13'h17A4: q=8'hE7;
	13'h17A5: q=8'hA8;
	13'h17A6: q=8'h86;
	13'h17A7: q=8'h55;
	13'h17A8: q=8'h97;
	13'h17A9: q=8'hEA;
	13'h17AA: q=8'h7E;
	13'h17AB: q=8'hE2;
	13'h17AC: q=8'h71;
	13'h17AD: q=8'hDD;
	13'h17AE: q=8'hBF;
	13'h17AF: q=8'hE6;
	13'h17B0: q=8'h0;
	13'h17B1: q=8'h8;
	13'h17B2: q=8'hA6;
	13'h17B3: q=8'h0;
	13'h17B4: q=8'hDF;
	13'h17B5: q=8'hC1;
	13'h17B6: q=8'hDE;
	13'h17B7: q=8'hBF;
	13'h17B8: q=8'hA7;
	13'h17B9: q=8'h0;
	13'h17BA: q=8'h8;
	13'h17BB: q=8'hDF;
	13'h17BC: q=8'hBF;
	13'h17BD: q=8'hDE;
	13'h17BE: q=8'hC1;
	13'h17BF: q=8'h5A;
	13'h17C0: q=8'h26;
	13'h17C1: q=8'hEF;
	13'h17C2: q=8'h39;
	13'h17C3: q=8'h1;
	13'h17C4: q=8'h7F;
	13'h17C5: q=8'h0;
	13'h17C6: q=8'hE8;
	13'h17C7: q=8'hBD;
	13'h17C8: q=8'hE3;
	13'h17C9: q=8'hEE;
	13'h17CA: q=8'hBD;
	13'h17CB: q=8'hFB;
	13'h17CC: q=8'hD4;
	13'h17CD: q=8'h20;
	13'h17CE: q=8'hDB;
	13'h17CF: q=8'hE;
	13'h17D0: q=8'h7C;
	13'h17D1: q=8'h0;
	13'h17D2: q=8'hF5;
	13'h17D3: q=8'h26;
	13'h17D4: q=8'h3;
	13'h17D5: q=8'h7C;
	13'h17D6: q=8'h0;
	13'h17D7: q=8'hF4;
	13'h17D8: q=8'hB6;
	13'h17D9: q=8'h0;
	13'h17DA: q=8'h0;
	13'h17DB: q=8'h7E;
	13'h17DC: q=8'hE1;
	13'h17DD: q=8'hC8;
	13'h17DE: q=8'h31;
	13'h17DF: q=8'h3B;
	13'h17E0: q=8'h0;
	13'h17E1: q=8'h0;
	13'h17E2: q=8'h3B;
	13'h17E3: q=8'h0;
	13'h17E4: q=8'h0;
	13'h17E5: q=8'h3B;
	13'h17E6: q=8'h0;
	13'h17E7: q=8'h0;
	13'h17E8: q=8'h3B;
	13'h17E9: q=8'h0;
	13'h17EA: q=8'h0;
	13'h17EB: q=8'h3B;
	13'h17EC: q=8'h0;
	13'h17ED: q=8'h0;
	13'h17EE: q=8'h3B;
	13'h17EF: q=8'h0;
	13'h17F0: q=8'h0;
	13'h17F1: q=8'h3B;
	13'h17F2: q=8'h0;
	13'h17F3: q=8'h0;
	13'h17F4: q=8'h7E;
	13'h17F5: q=8'hEC;
	13'h17F6: q=8'h2E;
	13'h17F7: q=8'h4F;
	13'h17F8: q=8'hC7;
	13'h17F9: q=8'h52;
	13'h17FA: q=8'h59;
	13'h17FB: q=8'hFF;
	13'h17FC: q=8'h4;
	13'h17FD: q=8'h5E;
	13'h17FE: q=8'hEC;
	13'h17FF: q=8'h2E;
	13'h1800: q=8'hF7;
	13'h1801: q=8'hC3;
	13'h1802: q=8'h0;
	13'h1803: q=8'h76;
	13'h1804: q=8'h0;
	13'h1805: q=8'h1;
	13'h1806: q=8'h10;
	13'h1807: q=8'h70;
	13'h1808: q=8'h84;
	13'h1809: q=8'h0;
	13'h180A: q=8'h1;
	13'h180B: q=8'h15;
	13'h180C: q=8'h1A;
	13'h180D: q=8'hB;
	13'h180E: q=8'h0;
	13'h180F: q=8'h80;
	13'h1810: q=8'h4D;
	13'h1811: q=8'h49;
	13'h1812: q=8'h43;
	13'h1813: q=8'h52;
	13'h1814: q=8'h4F;
	13'h1815: q=8'h43;
	13'h1816: q=8'h4F;
	13'h1817: q=8'h4C;
	13'h1818: q=8'h4F;
	13'h1819: q=8'h52;
	13'h181A: q=8'h20;
	13'h181B: q=8'h42;
	13'h181C: q=8'h41;
	13'h181D: q=8'h53;
	13'h181E: q=8'h49;
	13'h181F: q=8'h43;
	13'h1820: q=8'h20;
	13'h1821: q=8'h31;
	13'h1822: q=8'h2E;
	13'h1823: q=8'h30;
	13'h1824: q=8'hD;
	13'h1825: q=8'h43;
	13'h1826: q=8'h4F;
	13'h1827: q=8'h50;
	13'h1828: q=8'h59;
	13'h1829: q=8'h52;
	13'h182A: q=8'h49;
	13'h182B: q=8'h47;
	13'h182C: q=8'h48;
	13'h182D: q=8'h54;
	13'h182E: q=8'h20;
	13'h182F: q=8'h31;
	13'h1830: q=8'h39;
	13'h1831: q=8'h38;
	13'h1832: q=8'h32;
	13'h1833: q=8'h20;
	13'h1834: q=8'h4D;
	13'h1835: q=8'h49;
	13'h1836: q=8'h43;
	13'h1837: q=8'h52;
	13'h1838: q=8'h4F;
	13'h1839: q=8'h53;
	13'h183A: q=8'h4F;
	13'h183B: q=8'h46;
	13'h183C: q=8'h54;
	13'h183D: q=8'hD;
	13'h183E: q=8'h0;
	13'h183F: q=8'h7A;
	13'h1840: q=8'h42;
	13'h1841: q=8'h2B;
	13'h1842: q=8'h26;
	13'h1843: q=8'h1A;
	13'h1844: q=8'hB6;
	13'h1845: q=8'h42;
	13'h1846: q=8'h82;
	13'h1847: q=8'h88;
	13'h1848: q=8'hF;
	13'h1849: q=8'hB7;
	13'h184A: q=8'h42;
	13'h184B: q=8'h82;
	13'h184C: q=8'h8A;
	13'h184D: q=8'h80;
	13'h184E: q=8'hFE;
	13'h184F: q=8'h42;
	13'h1850: q=8'h80;
	13'h1851: q=8'hA7;
	13'h1852: q=8'h0;
	13'h1853: q=8'hC6;
	13'h1854: q=8'h16;
	13'h1855: q=8'h84;
	13'h1856: q=8'hF;
	13'h1857: q=8'h27;
	13'h1858: q=8'h2;
	13'h1859: q=8'hC6;
	13'h185A: q=8'h58;
	13'h185B: q=8'hF7;
	13'h185C: q=8'h42;
	13'h185D: q=8'h2B;
	13'h185E: q=8'hCE;
	13'h185F: q=8'h3;
	13'h1860: q=8'hFA;
	13'h1861: q=8'h9;
	13'h1862: q=8'h26;
	13'h1863: q=8'hFD;
	13'h1864: q=8'h39;
	13'h1865: q=8'hBD;
	13'h1866: q=8'h42;
	13'h1867: q=8'h85;
	13'h1868: q=8'h3C;
	13'h1869: q=8'h37;
	13'h186A: q=8'h8D;
	13'h186B: q=8'hD3;
	13'h186C: q=8'h8D;
	13'h186D: q=8'h15;
	13'h186E: q=8'h27;
	13'h186F: q=8'hFA;
	13'h1870: q=8'hC6;
	13'h1871: q=8'h60;
	13'h1872: q=8'hFE;
	13'h1873: q=8'h42;
	13'h1874: q=8'h80;
	13'h1875: q=8'hE7;
	13'h1876: q=8'h0;
	13'h1877: q=8'h20;
	13'h1878: q=8'h52;
	13'h1879: q=8'h4F;
	13'h187A: q=8'h8D;
	13'h187B: q=8'h54;
	13'h187C: q=8'h26;
	13'h187D: q=8'h5;
	13'h187E: q=8'h8D;
	13'h187F: q=8'h64;
	13'h1880: q=8'h4C;
	13'h1881: q=8'h27;
	13'h1882: q=8'h4A;
	13'h1883: q=8'hBD;
	13'h1884: q=8'h42;
	13'h1885: q=8'hA9;
	13'h1886: q=8'h3C;
	13'h1887: q=8'h37;
	13'h1888: q=8'h86;
	13'h1889: q=8'hFB;
	13'h188A: q=8'h8D;
	13'h188B: q=8'h44;
	13'h188C: q=8'h16;
	13'h188D: q=8'h27;
	13'h188E: q=8'h3;
	13'h188F: q=8'hF8;
	13'h1890: q=8'h42;
	13'h1891: q=8'h3B;
	13'h1892: q=8'hB7;
	13'h1893: q=8'h42;
	13'h1894: q=8'h3B;
	13'h1895: q=8'h5D;
	13'h1896: q=8'h27;
	13'h1897: q=8'h6;
	13'h1898: q=8'h8D;
	13'h1899: q=8'h42;
	13'h189A: q=8'h8D;
	13'h189B: q=8'h36;
	13'h189C: q=8'h26;
	13'h189D: q=8'h2A;
	13'h189E: q=8'hCE;
	13'h189F: q=8'h42;
	13'h18A0: q=8'h30;
	13'h18A1: q=8'h5F;
	13'h18A2: q=8'h5A;
	13'h18A3: q=8'hF7;
	13'h18A4: q=8'h42;
	13'h18A5: q=8'h39;
	13'h18A6: q=8'h59;
	13'h18A7: q=8'h24;
	13'h18A8: q=8'h1D;
	13'h18A9: q=8'h7C;
	13'h18AA: q=8'h42;
	13'h18AB: q=8'h39;
	13'h18AC: q=8'h8D;
	13'h18AD: q=8'h34;
	13'h18AE: q=8'h37;
	13'h18AF: q=8'h16;
	13'h18B0: q=8'h8;
	13'h18B1: q=8'hA8;
	13'h18B2: q=8'h0;
	13'h18B3: q=8'hA4;
	13'h18B4: q=8'h0;
	13'h18B5: q=8'hE7;
	13'h18B6: q=8'h0;
	13'h18B7: q=8'h33;
	13'h18B8: q=8'h4D;
	13'h18B9: q=8'hD;
	13'h18BA: q=8'h27;
	13'h18BB: q=8'hEA;
	13'h18BC: q=8'h36;
	13'h18BD: q=8'h8D;
	13'h18BE: q=8'h1D;
	13'h18BF: q=8'h8D;
	13'h18C0: q=8'h23;
	13'h18C1: q=8'hA1;
	13'h18C2: q=8'h0;
	13'h18C3: q=8'h32;
	13'h18C4: q=8'h26;
	13'h18C5: q=8'h24;
	13'h18C6: q=8'h4F;
	13'h18C7: q=8'h8C;
	13'h18C8: q=8'h86;
	13'h18C9: q=8'h3;
	13'h18CA: q=8'h4D;
	13'h18CB: q=8'h33;
	13'h18CC: q=8'h38;
	13'h18CD: q=8'h39;
	13'h18CE: q=8'h86;
	13'h18CF: q=8'h7F;
	13'h18D0: q=8'h97;
	13'h18D1: q=8'h2;
	13'h18D2: q=8'h96;
	13'h18D3: q=8'h3;
	13'h18D4: q=8'h43;
	13'h18D5: q=8'h84;
	13'h18D6: q=8'h2;
	13'h18D7: q=8'h27;
	13'h18D8: q=8'h2;
	13'h18D9: q=8'h86;
	13'h18DA: q=8'hFF;
	13'h18DB: q=8'h39;
	13'h18DC: q=8'hFE;
	13'h18DD: q=8'h42;
	13'h18DE: q=8'h1D;
	13'h18DF: q=8'h7E;
	13'h18E0: q=8'hF8;
	13'h18E1: q=8'h61;
	13'h18E2: q=8'hD7;
	13'h18E3: q=8'h2;
	13'h18E4: q=8'hB6;
	13'h18E5: q=8'hBF;
	13'h18E6: q=8'hFF;
	13'h18E7: q=8'h8A;
	13'h18E8: q=8'hC0;
	13'h18E9: q=8'h39;
	13'h18EA: q=8'hC6;
	13'h18EB: q=8'hF8;
	13'h18EC: q=8'hCB;
	13'h18ED: q=8'h8;
	13'h18EE: q=8'h44;
	13'h18EF: q=8'h24;
	13'h18F0: q=8'hFB;
	13'h18F1: q=8'hFB;
	13'h18F2: q=8'h42;
	13'h18F3: q=8'h39;
	13'h18F4: q=8'h86;
	13'h18F5: q=8'hFE;
	13'h18F6: q=8'h8D;
	13'h18F7: q=8'hD8;
	13'h18F8: q=8'hB7;
	13'h18F9: q=8'h42;
	13'h18FA: q=8'h3A;
	13'h18FB: q=8'hBD;
	13'h18FC: q=8'h42;
	13'h18FD: q=8'hAC;
	13'h18FE: q=8'h27;
	13'h18FF: q=8'h11;
	13'h1900: q=8'hCE;
	13'h1901: q=8'hF9;
	13'h1902: q=8'h7C;
	13'h1903: q=8'hC1;
	13'h1904: q=8'h20;
	13'h1905: q=8'h26;
	13'h1906: q=8'h27;
	13'h1907: q=8'hB6;
	13'h1908: q=8'h42;
	13'h1909: q=8'h82;
	13'h190A: q=8'h8B;
	13'h190B: q=8'h10;
	13'h190C: q=8'hB7;
	13'h190D: q=8'h42;
	13'h190E: q=8'h82;
	13'h190F: q=8'h20;
	13'h1910: q=8'hB5;
	13'h1911: q=8'h17;
	13'h1912: q=8'h27;
	13'h1913: q=8'h5;
	13'h1914: q=8'hC1;
	13'h1915: q=8'h1A;
	13'h1916: q=8'h23;
	13'h1917: q=8'h1B;
	13'h1918: q=8'h8C;
	13'h1919: q=8'hC6;
	13'h191A: q=8'h1D;
	13'h191B: q=8'hCE;
	13'h191C: q=8'hF9;
	13'h191D: q=8'h39;
	13'h191E: q=8'h8D;
	13'h191F: q=8'hAE;
	13'h1920: q=8'h27;
	13'h1921: q=8'hC;
	13'h1922: q=8'hCE;
	13'h1923: q=8'hF9;
	13'h1924: q=8'h4C;
	13'h1925: q=8'hC1;
	13'h1926: q=8'h20;
	13'h1927: q=8'h26;
	13'h1928: q=8'h5;
	13'h1929: q=8'h73;
	13'h192A: q=8'h42;
	13'h192B: q=8'h1C;
	13'h192C: q=8'h20;
	13'h192D: q=8'h98;
	13'h192E: q=8'h3A;
	13'h192F: q=8'hA6;
	13'h1930: q=8'h0;
	13'h1931: q=8'h20;
	13'h1932: q=8'h97;
	13'h1933: q=8'h8D;
	13'h1934: q=8'h99;
	13'h1935: q=8'hB8;
	13'h1936: q=8'h42;
	13'h1937: q=8'h1C;
	13'h1938: q=8'h26;
	13'h1939: q=8'h7;
	13'h193A: q=8'hB6;
	13'h193B: q=8'h42;
	13'h193C: q=8'h1C;
	13'h193D: q=8'h26;
	13'h193E: q=8'h7;
	13'h193F: q=8'hCA;
	13'h1940: q=8'h20;
	13'h1941: q=8'h17;
	13'h1942: q=8'h8A;
	13'h1943: q=8'h40;
	13'h1944: q=8'h20;
	13'h1945: q=8'h84;
	13'h1946: q=8'hCE;
	13'h1947: q=8'hF9;
	13'h1948: q=8'hAB;
	13'h1949: q=8'h3A;
	13'h194A: q=8'hA6;
	13'h194B: q=8'h0;
	13'h194C: q=8'h2A;
	13'h194D: q=8'hF6;
	13'h194E: q=8'hF6;
	13'h194F: q=8'h42;
	13'h1950: q=8'h82;
	13'h1951: q=8'hC4;
	13'h1952: q=8'h70;
	13'h1953: q=8'h1B;
	13'h1954: q=8'h20;
	13'h1955: q=8'hEE;
	13'h1956: q=8'h40;
	13'h1957: q=8'hD;
	13'h1958: q=8'h20;
	13'h1959: q=8'h30;
	13'h195A: q=8'h31;
	13'h195B: q=8'h32;
	13'h195C: q=8'h33;
	13'h195D: q=8'h34;
	13'h195E: q=8'h35;
	13'h195F: q=8'h36;
	13'h1960: q=8'h37;
	13'h1961: q=8'h38;
	13'h1962: q=8'h39;
	13'h1963: q=8'h3A;
	13'h1964: q=8'h3B;
	13'h1965: q=8'h2C;
	13'h1966: q=8'h2D;
	13'h1967: q=8'h2E;
	13'h1968: q=8'h2F;
	13'h1969: q=8'h13;
	13'h196A: q=8'hD;
	13'h196B: q=8'h20;
	13'h196C: q=8'h0;
	13'h196D: q=8'h21;
	13'h196E: q=8'h22;
	13'h196F: q=8'h23;
	13'h1970: q=8'h24;
	13'h1971: q=8'h25;
	13'h1972: q=8'h26;
	13'h1973: q=8'h27;
	13'h1974: q=8'h28;
	13'h1975: q=8'h29;
	13'h1976: q=8'h2A;
	13'h1977: q=8'h2B;
	13'h1978: q=8'h3C;
	13'h1979: q=8'h3D;
	13'h197A: q=8'h3E;
	13'h197B: q=8'h3F;
	13'h197C: q=8'h88;
	13'h197D: q=8'h8;
	13'h197E: q=8'hB3;
	13'h197F: q=8'hB2;
	13'h1980: q=8'h82;
	13'h1981: q=8'h9B;
	13'h1982: q=8'h90;
	13'h1983: q=8'h84;
	13'h1984: q=8'hA3;
	13'h1985: q=8'h8A;
	13'h1986: q=8'h81;
	13'h1987: q=8'h9E;
	13'h1988: q=8'hBC;
	13'h1989: q=8'hBA;
	13'h198A: q=8'hB9;
	13'h198B: q=8'hA5;
	13'h198C: q=8'hC7;
	13'h198D: q=8'h15;
	13'h198E: q=8'h9C;
	13'h198F: q=8'h9;
	13'h1990: q=8'h8C;
	13'h1991: q=8'h80;
	13'h1992: q=8'hB5;
	13'h1993: q=8'h5E;
	13'h1994: q=8'hB1;
	13'h1995: q=8'h8F;
	13'h1996: q=8'hA;
	13'h1997: q=8'h0;
	13'h1998: q=8'h0;
	13'h1999: q=8'h0;
	13'h199A: q=8'hD;
	13'h199B: q=8'h20;
	13'h199C: q=8'h0;
	13'h199D: q=8'h8E;
	13'h199E: q=8'h93;
	13'h199F: q=8'h98;
	13'h19A0: q=8'h97;
	13'h19A1: q=8'h96;
	13'h19A2: q=8'h94;
	13'h19A3: q=8'h95;
	13'h19A4: q=8'h9D;
	13'h19A5: q=8'h86;
	13'h19A6: q=8'h89;
	13'h19A7: q=8'h92;
	13'h19A8: q=8'hBB;
	13'h19A9: q=8'h91;
	13'h19AA: q=8'hB7;
	13'h19AB: q=8'hB6;
	13'h19AC: q=8'h89;
	13'h19AD: q=8'h80;
	13'h19AE: q=8'h82;
	13'h19AF: q=8'h87;
	13'h19B0: q=8'h8D;
	13'h19B1: q=8'h86;
	13'h19B2: q=8'h85;
	13'h19B3: q=8'h48;
	13'h19B4: q=8'h49;
	13'h19B5: q=8'h4A;
	13'h19B6: q=8'h4B;
	13'h19B7: q=8'h4C;
	13'h19B8: q=8'h4D;
	13'h19B9: q=8'h4E;
	13'h19BA: q=8'h4F;
	13'h19BB: q=8'h50;
	13'h19BC: q=8'h8F;
	13'h19BD: q=8'h8C;
	13'h19BE: q=8'h88;
	13'h19BF: q=8'h8B;
	13'h19C0: q=8'h55;
	13'h19C1: q=8'h81;
	13'h19C2: q=8'h8E;
	13'h19C3: q=8'h83;
	13'h19C4: q=8'h8A;
	13'h19C5: q=8'h84;
	13'h19C6: q=8'hBD;
	13'h19C7: q=8'h42;
	13'h19C8: q=8'h88;
	13'h19C9: q=8'h3C;
	13'h19CA: q=8'h37;
	13'h19CB: q=8'h36;
	13'h19CC: q=8'hD6;
	13'h19CD: q=8'hE8;
	13'h19CE: q=8'h27;
	13'h19CF: q=8'h4B;
	13'h19D0: q=8'h16;
	13'h19D1: q=8'h7;
	13'h19D2: q=8'h36;
	13'h19D3: q=8'hF;
	13'h19D4: q=8'h17;
	13'h19D5: q=8'hD6;
	13'h19D6: q=8'h3;
	13'h19D7: q=8'hC4;
	13'h19D8: q=8'h4;
	13'h19D9: q=8'h26;
	13'h19DA: q=8'hFA;
	13'h19DB: q=8'h8D;
	13'h19DC: q=8'h2D;
	13'h19DD: q=8'h5F;
	13'h19DE: q=8'h8D;
	13'h19DF: q=8'h2C;
	13'h19E0: q=8'hC6;
	13'h19E1: q=8'h8;
	13'h19E2: q=8'h37;
	13'h19E3: q=8'h5F;
	13'h19E4: q=8'h44;
	13'h19E5: q=8'h59;
	13'h19E6: q=8'h8D;
	13'h19E7: q=8'h24;
	13'h19E8: q=8'h33;
	13'h19E9: q=8'h5A;
	13'h19EA: q=8'h26;
	13'h19EB: q=8'hF6;
	13'h19EC: q=8'h8D;
	13'h19ED: q=8'h1C;
	13'h19EE: q=8'h32;
	13'h19EF: q=8'h6;
	13'h19F0: q=8'h32;
	13'h19F1: q=8'h81;
	13'h19F2: q=8'hD;
	13'h19F3: q=8'h27;
	13'h19F4: q=8'hB;
	13'h19F5: q=8'h7C;
	13'h19F6: q=8'h42;
	13'h19F7: q=8'h2A;
	13'h19F8: q=8'hF6;
	13'h19F9: q=8'h42;
	13'h19FA: q=8'h2A;
	13'h19FB: q=8'hF1;
	13'h19FC: q=8'h42;
	13'h19FD: q=8'h29;
	13'h19FE: q=8'h25;
	13'h19FF: q=8'h7;
	13'h1A00: q=8'h7F;
	13'h1A01: q=8'h42;
	13'h1A02: q=8'h2A;
	13'h1A03: q=8'h8D;
	13'h1A04: q=8'h10;
	13'h1A05: q=8'h8D;
	13'h1A06: q=8'hE;
	13'h1A07: q=8'h33;
	13'h1A08: q=8'h38;
	13'h1A09: q=8'h39;
	13'h1A0A: q=8'hC6;
	13'h1A0B: q=8'h1;
	13'h1A0C: q=8'hD7;
	13'h1A0D: q=8'h3;
	13'h1A0E: q=8'h8D;
	13'h1A0F: q=8'h0;
	13'h1A10: q=8'hFE;
	13'h1A11: q=8'h42;
	13'h1A12: q=8'h23;
	13'h1A13: q=8'h20;
	13'h1A14: q=8'h3;
	13'h1A15: q=8'hFE;
	13'h1A16: q=8'h42;
	13'h1A17: q=8'h25;
	13'h1A18: q=8'h7E;
	13'h1A19: q=8'hF8;
	13'h1A1A: q=8'h61;
	13'h1A1B: q=8'hFE;
	13'h1A1C: q=8'h42;
	13'h1A1D: q=8'h80;
	13'h1A1E: q=8'h81;
	13'h1A1F: q=8'h8;
	13'h1A20: q=8'h26;
	13'h1A21: q=8'hC;
	13'h1A22: q=8'h8C;
	13'h1A23: q=8'h40;
	13'h1A24: q=8'h0;
	13'h1A25: q=8'h27;
	13'h1A26: q=8'h50;
	13'h1A27: q=8'h86;
	13'h1A28: q=8'h60;
	13'h1A29: q=8'h9;
	13'h1A2A: q=8'hA7;
	13'h1A2B: q=8'h0;
	13'h1A2C: q=8'h20;
	13'h1A2D: q=8'h2E;
	13'h1A2E: q=8'h81;
	13'h1A2F: q=8'hD;
	13'h1A30: q=8'h26;
	13'h1A31: q=8'h14;
	13'h1A32: q=8'hFE;
	13'h1A33: q=8'h42;
	13'h1A34: q=8'h80;
	13'h1A35: q=8'h86;
	13'h1A36: q=8'h60;
	13'h1A37: q=8'hA7;
	13'h1A38: q=8'h0;
	13'h1A39: q=8'h8;
	13'h1A3A: q=8'hFF;
	13'h1A3B: q=8'h42;
	13'h1A3C: q=8'h80;
	13'h1A3D: q=8'hF6;
	13'h1A3E: q=8'h42;
	13'h1A3F: q=8'h81;
	13'h1A40: q=8'hC5;
	13'h1A41: q=8'h1F;
	13'h1A42: q=8'h26;
	13'h1A43: q=8'hF1;
	13'h1A44: q=8'h20;
	13'h1A45: q=8'h16;
	13'h1A46: q=8'h81;
	13'h1A47: q=8'h20;
	13'h1A48: q=8'h25;
	13'h1A49: q=8'h2D;
	13'h1A4A: q=8'h4D;
	13'h1A4B: q=8'h2B;
	13'h1A4C: q=8'hC;
	13'h1A4D: q=8'h81;
	13'h1A4E: q=8'h40;
	13'h1A4F: q=8'h25;
	13'h1A50: q=8'h6;
	13'h1A51: q=8'h81;
	13'h1A52: q=8'h60;
	13'h1A53: q=8'h25;
	13'h1A54: q=8'h4;
	13'h1A55: q=8'h84;
	13'h1A56: q=8'hDF;
	13'h1A57: q=8'h88;
	13'h1A58: q=8'h40;
	13'h1A59: q=8'hA7;
	13'h1A5A: q=8'h0;
	13'h1A5B: q=8'h8;
	13'h1A5C: q=8'hFF;
	13'h1A5D: q=8'h42;
	13'h1A5E: q=8'h80;
	13'h1A5F: q=8'h8C;
	13'h1A60: q=8'h42;
	13'h1A61: q=8'h0;
	13'h1A62: q=8'h26;
	13'h1A63: q=8'h13;
	13'h1A64: q=8'hCE;
	13'h1A65: q=8'h40;
	13'h1A66: q=8'h0;
	13'h1A67: q=8'hEC;
	13'h1A68: q=8'h20;
	13'h1A69: q=8'hED;
	13'h1A6A: q=8'h0;
	13'h1A6B: q=8'h8;
	13'h1A6C: q=8'h8;
	13'h1A6D: q=8'h8C;
	13'h1A6E: q=8'h41;
	13'h1A6F: q=8'hE0;
	13'h1A70: q=8'h26;
	13'h1A71: q=8'hF5;
	13'h1A72: q=8'hC6;
	13'h1A73: q=8'h60;
	13'h1A74: q=8'hBD;
	13'h1A75: q=8'hFB;
	13'h1A76: q=8'hD9;
	13'h1A77: q=8'h32;
	13'h1A78: q=8'h33;
	13'h1A79: q=8'h38;
	13'h1A7A: q=8'h39;
	13'h1A7B: q=8'hBD;
	13'h1A7C: q=8'h42;
	13'h1A7D: q=8'h8B;
	13'h1A7E: q=8'h3C;
	13'h1A7F: q=8'h37;
	13'h1A80: q=8'h36;
	13'h1A81: q=8'h96;
	13'h1A82: q=8'hE8;
	13'h1A83: q=8'h27;
	13'h1A84: q=8'h8;
	13'h1A85: q=8'hFE;
	13'h1A86: q=8'h42;
	13'h1A87: q=8'h27;
	13'h1A88: q=8'hFC;
	13'h1A89: q=8'h42;
	13'h1A8A: q=8'h29;
	13'h1A8B: q=8'h20;
	13'h1A8C: q=8'hA;
	13'h1A8D: q=8'hF6;
	13'h1A8E: q=8'h42;
	13'h1A8F: q=8'h81;
	13'h1A90: q=8'hC4;
	13'h1A91: q=8'h1F;
	13'h1A92: q=8'hCE;
	13'h1A93: q=8'h10;
	13'h1A94: q=8'h10;
	13'h1A95: q=8'h86;
	13'h1A96: q=8'h20;
	13'h1A97: q=8'hDF;
	13'h1A98: q=8'hE4;
	13'h1A99: q=8'hD7;
	13'h1A9A: q=8'hE6;
	13'h1A9B: q=8'h97;
	13'h1A9C: q=8'hE7;
	13'h1A9D: q=8'h32;
	13'h1A9E: q=8'h33;
	13'h1A9F: q=8'h38;
	13'h1AA0: q=8'h39;
	13'h1AA1: q=8'hBD;
	13'h1AA2: q=8'hFB;
	13'h1AA3: q=8'hD4;
	13'h1AA4: q=8'hBD;
	13'h1AA5: q=8'h42;
	13'h1AA6: q=8'h91;
	13'h1AA7: q=8'h7F;
	13'h1AA8: q=8'h42;
	13'h1AA9: q=8'h7F;
	13'h1AAA: q=8'hCE;
	13'h1AAB: q=8'h42;
	13'h1AAC: q=8'hB2;
	13'h1AAD: q=8'hC6;
	13'h1AAE: q=8'h1;
	13'h1AAF: q=8'hBD;
	13'h1AB0: q=8'hF8;
	13'h1AB1: q=8'h65;
	13'h1AB2: q=8'h7D;
	13'h1AB3: q=8'h0;
	13'h1AB4: q=8'hE9;
	13'h1AB5: q=8'h26;
	13'h1AB6: q=8'h4D;
	13'h1AB7: q=8'h7D;
	13'h1AB8: q=8'h0;
	13'h1AB9: q=8'hE8;
	13'h1ABA: q=8'h26;
	13'h1ABB: q=8'h44;
	13'h1ABC: q=8'h4D;
	13'h1ABD: q=8'h2A;
	13'h1ABE: q=8'h1E;
	13'h1ABF: q=8'h7D;
	13'h1AC0: q=8'h42;
	13'h1AC1: q=8'h3A;
	13'h1AC2: q=8'h27;
	13'h1AC3: q=8'h19;
	13'h1AC4: q=8'hBD;
	13'h1AC5: q=8'hE4;
	13'h1AC6: q=8'hB2;
	13'h1AC7: q=8'hA6;
	13'h1AC8: q=8'h0;
	13'h1AC9: q=8'h8;
	13'h1ACA: q=8'h3C;
	13'h1ACB: q=8'h36;
	13'h1ACC: q=8'h84;
	13'h1ACD: q=8'h7F;
	13'h1ACE: q=8'hDE;
	13'h1ACF: q=8'h89;
	13'h1AD0: q=8'h8D;
	13'h1AD1: q=8'h48;
	13'h1AD2: q=8'hDF;
	13'h1AD3: q=8'h89;
	13'h1AD4: q=8'h32;
	13'h1AD5: q=8'h38;
	13'h1AD6: q=8'h4D;
	13'h1AD7: q=8'h2A;
	13'h1AD8: q=8'hEE;
	13'h1AD9: q=8'hDE;
	13'h1ADA: q=8'h89;
	13'h1ADB: q=8'h20;
	13'h1ADC: q=8'hD2;
	13'h1ADD: q=8'h81;
	13'h1ADE: q=8'hC;
	13'h1ADF: q=8'h27;
	13'h1AE0: q=8'hC0;
	13'h1AE1: q=8'h81;
	13'h1AE2: q=8'h8;
	13'h1AE3: q=8'h26;
	13'h1AE4: q=8'h8;
	13'h1AE5: q=8'h5A;
	13'h1AE6: q=8'h27;
	13'h1AE7: q=8'hBF;
	13'h1AE8: q=8'h9;
	13'h1AE9: q=8'h8D;
	13'h1AEA: q=8'h37;
	13'h1AEB: q=8'h20;
	13'h1AEC: q=8'hC2;
	13'h1AED: q=8'h81;
	13'h1AEE: q=8'h15;
	13'h1AEF: q=8'h26;
	13'h1AF0: q=8'hA;
	13'h1AF1: q=8'h5A;
	13'h1AF2: q=8'h27;
	13'h1AF3: q=8'hB3;
	13'h1AF4: q=8'h86;
	13'h1AF5: q=8'h8;
	13'h1AF6: q=8'hBD;
	13'h1AF7: q=8'hF9;
	13'h1AF8: q=8'hC6;
	13'h1AF9: q=8'h20;
	13'h1AFA: q=8'hF6;
	13'h1AFB: q=8'h81;
	13'h1AFC: q=8'h3;
	13'h1AFD: q=8'hD;
	13'h1AFE: q=8'h27;
	13'h1AFF: q=8'h5;
	13'h1B00: q=8'h81;
	13'h1B01: q=8'hD;
	13'h1B02: q=8'h26;
	13'h1B03: q=8'hE;
	13'h1B04: q=8'h4F;
	13'h1B05: q=8'h7;
	13'h1B06: q=8'h36;
	13'h1B07: q=8'hBD;
	13'h1B08: q=8'hE7;
	13'h1B09: q=8'h66;
	13'h1B0A: q=8'h6F;
	13'h1B0B: q=8'h0;
	13'h1B0C: q=8'hCE;
	13'h1B0D: q=8'h42;
	13'h1B0E: q=8'hB1;
	13'h1B0F: q=8'h32;
	13'h1B10: q=8'h6;
	13'h1B11: q=8'h39;
	13'h1B12: q=8'h81;
	13'h1B13: q=8'h20;
	13'h1B14: q=8'h25;
	13'h1B15: q=8'h99;
	13'h1B16: q=8'h8D;
	13'h1B17: q=8'h2;
	13'h1B18: q=8'h20;
	13'h1B19: q=8'h95;
	13'h1B1A: q=8'hC1;
	13'h1B1B: q=8'h80;
	13'h1B1C: q=8'h24;
	13'h1B1D: q=8'hF3;
	13'h1B1E: q=8'hA7;
	13'h1B1F: q=8'h0;
	13'h1B20: q=8'h8;
	13'h1B21: q=8'h5C;
	13'h1B22: q=8'h7E;
	13'h1B23: q=8'hF9;
	13'h1B24: q=8'hC6;
	13'h1B25: q=8'h8D;
	13'h1B26: q=8'h43;
	13'h1B27: q=8'h3C;
	13'h1B28: q=8'hBD;
	13'h1B29: q=8'hEF;
	13'h1B2A: q=8'h47;
	13'h1B2B: q=8'h38;
	13'h1B2C: q=8'hC1;
	13'h1B2D: q=8'h8;
	13'h1B2E: q=8'h22;
	13'h1B2F: q=8'h37;
	13'h1B30: q=8'h5A;
	13'h1B31: q=8'h2B;
	13'h1B32: q=8'h5;
	13'h1B33: q=8'h86;
	13'h1B34: q=8'h10;
	13'h1B35: q=8'h3D;
	13'h1B36: q=8'h20;
	13'h1B37: q=8'h8;
	13'h1B38: q=8'hE6;
	13'h1B39: q=8'h0;
	13'h1B3A: q=8'h2A;
	13'h1B3B: q=8'h3;
	13'h1B3C: q=8'hC4;
	13'h1B3D: q=8'h70;
	13'h1B3E: q=8'h21;
	13'h1B3F: q=8'h5F;
	13'h1B40: q=8'hD7;
	13'h1B41: q=8'h82;
	13'h1B42: q=8'h8D;
	13'h1B43: q=8'h70;
	13'h1B44: q=8'hA6;
	13'h1B45: q=8'h0;
	13'h1B46: q=8'h2B;
	13'h1B47: q=8'h1;
	13'h1B48: q=8'h4F;
	13'h1B49: q=8'h84;
	13'h1B4A: q=8'hF;
	13'h1B4B: q=8'hBA;
	13'h1B4C: q=8'h42;
	13'h1B4D: q=8'h3C;
	13'h1B4E: q=8'h9A;
	13'h1B4F: q=8'h82;
	13'h1B50: q=8'h8A;
	13'h1B51: q=8'h80;
	13'h1B52: q=8'hA7;
	13'h1B53: q=8'h0;
	13'h1B54: q=8'h39;
	13'h1B55: q=8'h8D;
	13'h1B56: q=8'h13;
	13'h1B57: q=8'h8D;
	13'h1B58: q=8'h5B;
	13'h1B59: q=8'h4F;
	13'h1B5A: q=8'hE6;
	13'h1B5B: q=8'h0;
	13'h1B5C: q=8'h2A;
	13'h1B5D: q=8'hF2;
	13'h1B5E: q=8'h73;
	13'h1B5F: q=8'h42;
	13'h1B60: q=8'h3C;
	13'h1B61: q=8'hF4;
	13'h1B62: q=8'h42;
	13'h1B63: q=8'h3C;
	13'h1B64: q=8'hE7;
	13'h1B65: q=8'h0;
	13'h1B66: q=8'h39;
	13'h1B67: q=8'h7E;
	13'h1B68: q=8'hEC;
	13'h1B69: q=8'h2E;
	13'h1B6A: q=8'hBD;
	13'h1B6B: q=8'hEA;
	13'h1B6C: q=8'h2C;
	13'h1B6D: q=8'hBD;
	13'h1B6E: q=8'hEF;
	13'h1B6F: q=8'hD;
	13'h1B70: q=8'hC1;
	13'h1B71: q=8'h3F;
	13'h1B72: q=8'h22;
	13'h1B73: q=8'hF3;
	13'h1B74: q=8'h37;
	13'h1B75: q=8'hBD;
	13'h1B76: q=8'hEF;
	13'h1B77: q=8'h47;
	13'h1B78: q=8'hC1;
	13'h1B79: q=8'h1F;
	13'h1B7A: q=8'h22;
	13'h1B7B: q=8'hEB;
	13'h1B7C: q=8'h37;
	13'h1B7D: q=8'h54;
	13'h1B7E: q=8'h86;
	13'h1B7F: q=8'h20;
	13'h1B80: q=8'h3D;
	13'h1B81: q=8'hC3;
	13'h1B82: q=8'h40;
	13'h1B83: q=8'h0;
	13'h1B84: q=8'h37;
	13'h1B85: q=8'h36;
	13'h1B86: q=8'h30;
	13'h1B87: q=8'hE6;
	13'h1B88: q=8'h3;
	13'h1B89: q=8'h54;
	13'h1B8A: q=8'h38;
	13'h1B8B: q=8'h3A;
	13'h1B8C: q=8'h32;
	13'h1B8D: q=8'h33;
	13'h1B8E: q=8'h84;
	13'h1B8F: q=8'h1;
	13'h1B90: q=8'h56;
	13'h1B91: q=8'h49;
	13'h1B92: q=8'hC6;
	13'h1B93: q=8'h10;
	13'h1B94: q=8'h54;
	13'h1B95: q=8'h4A;
	13'h1B96: q=8'h2A;
	13'h1B97: q=8'hFC;
	13'h1B98: q=8'hF7;
	13'h1B99: q=8'h42;
	13'h1B9A: q=8'h3C;
	13'h1B9B: q=8'h39;
	13'h1B9C: q=8'h8D;
	13'h1B9D: q=8'hCF;
	13'h1B9E: q=8'hC6;
	13'h1B9F: q=8'hFF;
	13'h1BA0: q=8'hA6;
	13'h1BA1: q=8'h0;
	13'h1BA2: q=8'h2A;
	13'h1BA3: q=8'hE;
	13'h1BA4: q=8'hB4;
	13'h1BA5: q=8'h42;
	13'h1BA6: q=8'h3C;
	13'h1BA7: q=8'h27;
	13'h1BA8: q=8'h8;
	13'h1BA9: q=8'hE6;
	13'h1BAA: q=8'h0;
	13'h1BAB: q=8'h54;
	13'h1BAC: q=8'h54;
	13'h1BAD: q=8'h54;
	13'h1BAE: q=8'h54;
	13'h1BAF: q=8'hC4;
	13'h1BB0: q=8'h7;
	13'h1BB1: q=8'h5C;
	13'h1BB2: q=8'h8D;
	13'h1BB3: q=8'h3;
	13'h1BB4: q=8'h7E;
	13'h1BB5: q=8'hEA;
	13'h1BB6: q=8'h29;
	13'h1BB7: q=8'h4F;
	13'h1BB8: q=8'h5D;
	13'h1BB9: q=8'h2A;
	13'h1BBA: q=8'h1;
	13'h1BBB: q=8'h43;
	13'h1BBC: q=8'h7E;
	13'h1BBD: q=8'hEC;
	13'h1BBE: q=8'hE3;
	13'h1BBF: q=8'h27;
	13'h1BC0: q=8'h13;
	13'h1BC1: q=8'hBD;
	13'h1BC2: q=8'hEF;
	13'h1BC3: q=8'hD;
	13'h1BC4: q=8'hC1;
	13'h1BC5: q=8'h8;
	13'h1BC6: q=8'h22;
	13'h1BC7: q=8'h1D;
	13'h1BC8: q=8'h5D;
	13'h1BC9: q=8'h27;
	13'h1BCA: q=8'h6;
	13'h1BCB: q=8'h5A;
	13'h1BCC: q=8'h86;
	13'h1BCD: q=8'h10;
	13'h1BCE: q=8'h3D;
	13'h1BCF: q=8'hCA;
	13'h1BD0: q=8'hF;
	13'h1BD1: q=8'hCA;
	13'h1BD2: q=8'h80;
	13'h1BD3: q=8'h8C;
	13'h1BD4: q=8'hC6;
	13'h1BD5: q=8'h60;
	13'h1BD6: q=8'hCE;
	13'h1BD7: q=8'h40;
	13'h1BD8: q=8'h0;
	13'h1BD9: q=8'hFF;
	13'h1BDA: q=8'h42;
	13'h1BDB: q=8'h80;
	13'h1BDC: q=8'hE7;
	13'h1BDD: q=8'h0;
	13'h1BDE: q=8'h8;
	13'h1BDF: q=8'h8C;
	13'h1BE0: q=8'h42;
	13'h1BE1: q=8'h0;
	13'h1BE2: q=8'h26;
	13'h1BE3: q=8'hF8;
	13'h1BE4: q=8'h39;
	13'h1BE5: q=8'h8D;
	13'h1BE6: q=8'hED;
	13'h1BE7: q=8'hCE;
	13'h1BE8: q=8'hF8;
	13'h1BE9: q=8'h33;
	13'h1BEA: q=8'h7E;
	13'h1BEB: q=8'hE7;
	13'h1BEC: q=8'hA8;
	13'h1BED: q=8'hB6;
	13'h1BEE: q=8'h42;
	13'h1BEF: q=8'h7F;
	13'h1BF0: q=8'h26;
	13'h1BF1: q=8'h3;
	13'h1BF2: q=8'hBD;
	13'h1BF3: q=8'hF8;
	13'h1BF4: q=8'h83;
	13'h1BF5: q=8'h7F;
	13'h1BF6: q=8'h42;
	13'h1BF7: q=8'h7F;
	13'h1BF8: q=8'h97;
	13'h1BF9: q=8'hCD;
	13'h1BFA: q=8'h27;
	13'h1BFB: q=8'h3;
	13'h1BFC: q=8'h7E;
	13'h1BFD: q=8'hEE;
	13'h1BFE: q=8'h91;
	13'h1BFF: q=8'h97;
	13'h1C00: q=8'hD0;
	13'h1C01: q=8'h7E;
	13'h1C02: q=8'hEE;
	13'h1C03: q=8'h9D;
	13'h1C04: q=8'h27;
	13'h1C05: q=8'h6;
	13'h1C06: q=8'hBD;
	13'h1C07: q=8'hEF;
	13'h1C08: q=8'h4C;
	13'h1C09: q=8'hFF;
	13'h1C0A: q=8'h42;
	13'h1C0B: q=8'h1F;
	13'h1C0C: q=8'hFE;
	13'h1C0D: q=8'h42;
	13'h1C0E: q=8'h1F;
	13'h1C0F: q=8'h6E;
	13'h1C10: q=8'h0;
	13'h1C11: q=8'hDE;
	13'h1C12: q=8'h99;
	13'h1C13: q=8'h3C;
	13'h1C14: q=8'hBD;
	13'h1C15: q=8'hEB;
	13'h1C16: q=8'h1B;
	13'h1C17: q=8'hBD;
	13'h1C18: q=8'hEA;
	13'h1C19: q=8'h29;
	13'h1C1A: q=8'hDF;
	13'h1C1B: q=8'h89;
	13'h1C1C: q=8'h38;
	13'h1C1D: q=8'hDC;
	13'h1C1E: q=8'h89;
	13'h1C1F: q=8'h9C;
	13'h1C20: q=8'h99;
	13'h1C21: q=8'h27;
	13'h1C22: q=8'h3;
	13'h1C23: q=8'h7E;
	13'h1C24: q=8'hEC;
	13'h1C25: q=8'h2E;
	13'h1C26: q=8'h7E;
	13'h1C27: q=8'hEC;
	13'h1C28: q=8'hE3;
	13'h1C29: q=8'hBD;
	13'h1C2A: q=8'hEB;
	13'h1C2B: q=8'hBA;
	13'h1C2C: q=8'h83;
	13'h1C2D: q=8'h1;
	13'h1C2E: q=8'hFF;
	13'h1C2F: q=8'h23;
	13'h1C30: q=8'h3;
	13'h1C31: q=8'h7E;
	13'h1C32: q=8'hEC;
	13'h1C33: q=8'h2E;
	13'h1C34: q=8'hC3;
	13'h1C35: q=8'h41;
	13'h1C36: q=8'hFF;
	13'h1C37: q=8'hFD;
	13'h1C38: q=8'h42;
	13'h1C39: q=8'h80;
	13'h1C3A: q=8'h39;
	13'h1C3B: q=8'hDE;
	13'h1C3C: q=8'h93;
	13'h1C3D: q=8'hFF;
	13'h1C3E: q=8'h42;
	13'h1C3F: q=8'h6F;
	13'h1C40: q=8'hDE;
	13'h1C41: q=8'h95;
	13'h1C42: q=8'hFF;
	13'h1C43: q=8'h42;
	13'h1C44: q=8'h71;
	13'h1C45: q=8'h5F;
	13'h1C46: q=8'h81;
	13'h1C47: q=8'hA9;
	13'h1C48: q=8'h26;
	13'h1C49: q=8'h5;
	13'h1C4A: q=8'hBD;
	13'h1C4B: q=8'hFD;
	13'h1C4C: q=8'hDB;
	13'h1C4D: q=8'hC6;
	13'h1C4E: q=8'h4;
	13'h1C4F: q=8'hF7;
	13'h1C50: q=8'h42;
	13'h1C51: q=8'h67;
	13'h1C52: q=8'hFC;
	13'h1C53: q=8'h42;
	13'h1C54: q=8'h71;
	13'h1C55: q=8'hB3;
	13'h1C56: q=8'h42;
	13'h1C57: q=8'h6F;
	13'h1C58: q=8'hFD;
	13'h1C59: q=8'h42;
	13'h1C5A: q=8'h6C;
	13'h1C5B: q=8'h8D;
	13'h1C5C: q=8'h2E;
	13'h1C5D: q=8'hFE;
	13'h1C5E: q=8'h42;
	13'h1C5F: q=8'h6F;
	13'h1C60: q=8'hFF;
	13'h1C61: q=8'h42;
	13'h1C62: q=8'h78;
	13'h1C63: q=8'h86;
	13'h1C64: q=8'hFF;
	13'h1C65: q=8'hB7;
	13'h1C66: q=8'h42;
	13'h1C67: q=8'h76;
	13'h1C68: q=8'hFC;
	13'h1C69: q=8'h42;
	13'h1C6A: q=8'h71;
	13'h1C6B: q=8'hB3;
	13'h1C6C: q=8'h42;
	13'h1C6D: q=8'h78;
	13'h1C6E: q=8'h23;
	13'h1C6F: q=8'hE;
	13'h1C70: q=8'h4D;
	13'h1C71: q=8'h26;
	13'h1C72: q=8'h7;
	13'h1C73: q=8'hC1;
	13'h1C74: q=8'hFF;
	13'h1C75: q=8'h27;
	13'h1C76: q=8'h3;
	13'h1C77: q=8'hF7;
	13'h1C78: q=8'h42;
	13'h1C79: q=8'h76;
	13'h1C7A: q=8'h8D;
	13'h1C7B: q=8'h44;
	13'h1C7C: q=8'h20;
	13'h1C7D: q=8'hE2;
	13'h1C7E: q=8'h70;
	13'h1C7F: q=8'h42;
	13'h1C80: q=8'h75;
	13'h1C81: q=8'h7F;
	13'h1C82: q=8'h42;
	13'h1C83: q=8'h76;
	13'h1C84: q=8'h8D;
	13'h1C85: q=8'h3A;
	13'h1C86: q=8'h86;
	13'h1C87: q=8'h1;
	13'h1C88: q=8'h97;
	13'h1C89: q=8'h3;
	13'h1C8A: q=8'h39;
	13'h1C8B: q=8'hBD;
	13'h1C8C: q=8'hFD;
	13'h1C8D: q=8'h29;
	13'h1C8E: q=8'hCE;
	13'h1C8F: q=8'h42;
	13'h1C90: q=8'h5F;
	13'h1C91: q=8'hFF;
	13'h1C92: q=8'h42;
	13'h1C93: q=8'h78;
	13'h1C94: q=8'hDF;
	13'h1C95: q=8'hBF;
	13'h1C96: q=8'h6F;
	13'h1C97: q=8'h9;
	13'h1C98: q=8'h6F;
	13'h1C99: q=8'hA;
	13'h1C9A: q=8'hCE;
	13'h1C9B: q=8'h42;
	13'h1C9C: q=8'h57;
	13'h1C9D: q=8'hC6;
	13'h1C9E: q=8'h8;
	13'h1C9F: q=8'hBD;
	13'h1CA0: q=8'hF7;
	13'h1CA1: q=8'hB2;
	13'h1CA2: q=8'h7F;
	13'h1CA3: q=8'h42;
	13'h1CA4: q=8'h75;
	13'h1CA5: q=8'h86;
	13'h1CA6: q=8'hF;
	13'h1CA7: q=8'hB7;
	13'h1CA8: q=8'h42;
	13'h1CA9: q=8'h76;
	13'h1CAA: q=8'h8D;
	13'h1CAB: q=8'hB;
	13'h1CAC: q=8'h8D;
	13'h1CAD: q=8'h12;
	13'h1CAE: q=8'h7C;
	13'h1CAF: q=8'h42;
	13'h1CB0: q=8'h75;
	13'h1CB1: q=8'hCE;
	13'h1CB2: q=8'h0;
	13'h1CB3: q=8'h0;
	13'h1CB4: q=8'hBD;
	13'h1CB5: q=8'hF8;
	13'h1CB6: q=8'h61;
	13'h1CB7: q=8'hFE;
	13'h1CB8: q=8'h42;
	13'h1CB9: q=8'h2F;
	13'h1CBA: q=8'h8D;
	13'h1CBB: q=8'h45;
	13'h1CBC: q=8'h9;
	13'h1CBD: q=8'h26;
	13'h1CBE: q=8'hFB;
	13'h1CBF: q=8'h39;
	13'h1CC0: q=8'h1;
	13'h1CC1: q=8'hF;
	13'h1CC2: q=8'hF6;
	13'h1CC3: q=8'h42;
	13'h1CC4: q=8'h76;
	13'h1CC5: q=8'hF7;
	13'h1CC6: q=8'h42;
	13'h1CC7: q=8'h7B;
	13'h1CC8: q=8'hB6;
	13'h1CC9: q=8'h42;
	13'h1CCA: q=8'h76;
	13'h1CCB: q=8'h27;
	13'h1CCC: q=8'h9;
	13'h1CCD: q=8'hFE;
	13'h1CCE: q=8'h42;
	13'h1CCF: q=8'h78;
	13'h1CD0: q=8'hAB;
	13'h1CD1: q=8'h0;
	13'h1CD2: q=8'h8;
	13'h1CD3: q=8'h5A;
	13'h1CD4: q=8'h26;
	13'h1CD5: q=8'hFA;
	13'h1CD6: q=8'hBB;
	13'h1CD7: q=8'h42;
	13'h1CD8: q=8'h75;
	13'h1CD9: q=8'hB7;
	13'h1CDA: q=8'h42;
	13'h1CDB: q=8'h7A;
	13'h1CDC: q=8'hFE;
	13'h1CDD: q=8'h42;
	13'h1CDE: q=8'h78;
	13'h1CDF: q=8'h8D;
	13'h1CE0: q=8'h20;
	13'h1CE1: q=8'h86;
	13'h1CE2: q=8'h3C;
	13'h1CE3: q=8'h8D;
	13'h1CE4: q=8'h1E;
	13'h1CE5: q=8'hB6;
	13'h1CE6: q=8'h42;
	13'h1CE7: q=8'h75;
	13'h1CE8: q=8'h8D;
	13'h1CE9: q=8'h19;
	13'h1CEA: q=8'hB6;
	13'h1CEB: q=8'h42;
	13'h1CEC: q=8'h76;
	13'h1CED: q=8'h8D;
	13'h1CEE: q=8'h14;
	13'h1CEF: q=8'h4D;
	13'h1CF0: q=8'h27;
	13'h1CF1: q=8'hA;
	13'h1CF2: q=8'hA6;
	13'h1CF3: q=8'h0;
	13'h1CF4: q=8'h8;
	13'h1CF5: q=8'h8D;
	13'h1CF6: q=8'hC;
	13'h1CF7: q=8'h7A;
	13'h1CF8: q=8'h42;
	13'h1CF9: q=8'h7B;
	13'h1CFA: q=8'h26;
	13'h1CFB: q=8'hF6;
	13'h1CFC: q=8'hB6;
	13'h1CFD: q=8'h42;
	13'h1CFE: q=8'h7A;
	13'h1CFF: q=8'h8D;
	13'h1D00: q=8'h2;
	13'h1D01: q=8'h86;
	13'h1D02: q=8'h55;
	13'h1D03: q=8'h3C;
	13'h1D04: q=8'h36;
	13'h1D05: q=8'h36;
	13'h1D06: q=8'hC6;
	13'h1D07: q=8'h8;
	13'h1D08: q=8'h30;
	13'h1D09: q=8'h64;
	13'h1D0A: q=8'h0;
	13'h1D0B: q=8'hCE;
	13'h1D0C: q=8'h0;
	13'h1D0D: q=8'h20;
	13'h1D0E: q=8'h25;
	13'h1D0F: q=8'h3;
	13'h1D10: q=8'hCE;
	13'h1D11: q=8'h0;
	13'h1D12: q=8'h40;
	13'h1D13: q=8'h3C;
	13'h1D14: q=8'h86;
	13'h1D15: q=8'h1;
	13'h1D16: q=8'h97;
	13'h1D17: q=8'h3;
	13'h1D18: q=8'h9;
	13'h1D19: q=8'h26;
	13'h1D1A: q=8'hFD;
	13'h1D1B: q=8'h4F;
	13'h1D1C: q=8'h97;
	13'h1D1D: q=8'h3;
	13'h1D1E: q=8'h38;
	13'h1D1F: q=8'h9;
	13'h1D20: q=8'h26;
	13'h1D21: q=8'hFD;
	13'h1D22: q=8'h5A;
	13'h1D23: q=8'h26;
	13'h1D24: q=8'hE3;
	13'h1D25: q=8'h32;
	13'h1D26: q=8'h32;
	13'h1D27: q=8'h38;
	13'h1D28: q=8'h39;
	13'h1D29: q=8'h8D;
	13'h1D2A: q=8'h8;
	13'h1D2B: q=8'hBD;
	13'h1D2C: q=8'h0;
	13'h1D2D: q=8'hF3;
	13'h1D2E: q=8'h27;
	13'h1D2F: q=8'hF8;
	13'h1D30: q=8'h7E;
	13'h1D31: q=8'hEA;
	13'h1D32: q=8'h3C;
	13'h1D33: q=8'hCE;
	13'h1D34: q=8'h42;
	13'h1D35: q=8'h56;
	13'h1D36: q=8'h6F;
	13'h1D37: q=8'h0;
	13'h1D38: q=8'h86;
	13'h1D39: q=8'h20;
	13'h1D3A: q=8'h8;
	13'h1D3B: q=8'hA7;
	13'h1D3C: q=8'h0;
	13'h1D3D: q=8'h8C;
	13'h1D3E: q=8'h42;
	13'h1D3F: q=8'h5F;
	13'h1D40: q=8'h26;
	13'h1D41: q=8'hF8;
	13'h1D42: q=8'hBD;
	13'h1D43: q=8'h0;
	13'h1D44: q=8'hF3;
	13'h1D45: q=8'h27;
	13'h1D46: q=8'hE1;
	13'h1D47: q=8'hBD;
	13'h1D48: q=8'hE9;
	13'h1D49: q=8'h1A;
	13'h1D4A: q=8'hBD;
	13'h1D4B: q=8'hEE;
	13'h1D4C: q=8'h53;
	13'h1D4D: q=8'hF7;
	13'h1D4E: q=8'h42;
	13'h1D4F: q=8'h56;
	13'h1D50: q=8'h27;
	13'h1D51: q=8'hD6;
	13'h1D52: q=8'h37;
	13'h1D53: q=8'hCC;
	13'h1D54: q=8'h42;
	13'h1D55: q=8'h57;
	13'h1D56: q=8'hDD;
	13'h1D57: q=8'hBF;
	13'h1D58: q=8'h33;
	13'h1D59: q=8'h7E;
	13'h1D5A: q=8'hF7;
	13'h1D5B: q=8'hB2;
	13'h1D5C: q=8'h81;
	13'h1D5D: q=8'hA9;
	13'h1D5E: q=8'h26;
	13'h1D5F: q=8'h3;
	13'h1D60: q=8'h7E;
	13'h1D61: q=8'hFD;
	13'h1D62: q=8'hB1;
	13'h1D63: q=8'h81;
	13'h1D64: q=8'h4D;
	13'h1D65: q=8'h26;
	13'h1D66: q=8'h3;
	13'h1D67: q=8'h7E;
	13'h1D68: q=8'hFE;
	13'h1D69: q=8'h6;
	13'h1D6A: q=8'h4F;
	13'h1D6B: q=8'h8D;
	13'h1D6C: q=8'h22;
	13'h1D6D: q=8'hBD;
	13'h1D6E: q=8'hE3;
	13'h1D6F: q=8'hCF;
	13'h1D70: q=8'h73;
	13'h1D71: q=8'h42;
	13'h1D72: q=8'h6E;
	13'h1D73: q=8'hFC;
	13'h1D74: q=8'h42;
	13'h1D75: q=8'h6C;
	13'h1D76: q=8'hD3;
	13'h1D77: q=8'h93;
	13'h1D78: q=8'hBD;
	13'h1D79: q=8'hE2;
	13'h1D7A: q=8'h1E;
	13'h1D7B: q=8'hDE;
	13'h1D7C: q=8'h93;
	13'h1D7D: q=8'hFF;
	13'h1D7E: q=8'h42;
	13'h1D7F: q=8'h78;
	13'h1D80: q=8'h8D;
	13'h1D81: q=8'h4E;
	13'h1D82: q=8'h2A;
	13'h1D83: q=8'hF9;
	13'h1D84: q=8'hDF;
	13'h1D85: q=8'h95;
	13'h1D86: q=8'hCE;
	13'h1D87: q=8'hE1;
	13'h1D88: q=8'hBB;
	13'h1D89: q=8'hBD;
	13'h1D8A: q=8'hE7;
	13'h1D8B: q=8'hA8;
	13'h1D8C: q=8'h7E;
	13'h1D8D: q=8'hE2;
	13'h1D8E: q=8'hEB;
	13'h1D8F: q=8'h36;
	13'h1D90: q=8'h8D;
	13'h1D91: q=8'h10;
	13'h1D92: q=8'h32;
	13'h1D93: q=8'h7D;
	13'h1D94: q=8'h42;
	13'h1D95: q=8'h74;
	13'h1D96: q=8'h26;
	13'h1D97: q=8'h37;
	13'h1D98: q=8'hB1;
	13'h1D99: q=8'h42;
	13'h1D9A: q=8'h67;
	13'h1D9B: q=8'h27;
	13'h1D9C: q=8'h32;
	13'h1D9D: q=8'hC6;
	13'h1D9E: q=8'h24;
	13'h1D9F: q=8'h7E;
	13'h1DA0: q=8'hE2;
	13'h1DA1: q=8'h38;
	13'h1DA2: q=8'h8D;
	13'h1DA3: q=8'h8F;
	13'h1DA4: q=8'hBD;
	13'h1DA5: q=8'hFE;
	13'h1DA6: q=8'h37;
	13'h1DA7: q=8'h26;
	13'h1DA8: q=8'h3;
	13'h1DA9: q=8'h7E;
	13'h1DAA: q=8'hFF;
	13'h1DAB: q=8'h4E;
	13'h1DAC: q=8'hC6;
	13'h1DAD: q=8'h22;
	13'h1DAE: q=8'h7E;
	13'h1DAF: q=8'hE2;
	13'h1DB0: q=8'h38;
	13'h1DB1: q=8'h8D;
	13'h1DB2: q=8'h28;
	13'h1DB3: q=8'h86;
	13'h1DB4: q=8'h4;
	13'h1DB5: q=8'h8D;
	13'h1DB6: q=8'hD8;
	13'h1DB7: q=8'hFC;
	13'h1DB8: q=8'h42;
	13'h1DB9: q=8'h71;
	13'h1DBA: q=8'hB3;
	13'h1DBB: q=8'h42;
	13'h1DBC: q=8'h6F;
	13'h1DBD: q=8'hB3;
	13'h1DBE: q=8'h42;
	13'h1DBF: q=8'h6C;
	13'h1DC0: q=8'h24;
	13'h1DC1: q=8'h3;
	13'h1DC2: q=8'h7E;
	13'h1DC3: q=8'hE2;
	13'h1DC4: q=8'h36;
	13'h1DC5: q=8'hFE;
	13'h1DC6: q=8'h42;
	13'h1DC7: q=8'h6F;
	13'h1DC8: q=8'hFF;
	13'h1DC9: q=8'h42;
	13'h1DCA: q=8'h78;
	13'h1DCB: q=8'h8D;
	13'h1DCC: q=8'h3;
	13'h1DCD: q=8'h2A;
	13'h1DCE: q=8'hF9;
	13'h1DCF: q=8'h39;
	13'h1DD0: q=8'hBD;
	13'h1DD1: q=8'hFE;
	13'h1DD2: q=8'hB6;
	13'h1DD3: q=8'h26;
	13'h1DD4: q=8'hD7;
	13'h1DD5: q=8'hB6;
	13'h1DD6: q=8'h42;
	13'h1DD7: q=8'h75;
	13'h1DD8: q=8'h27;
	13'h1DD9: q=8'hD2;
	13'h1DDA: q=8'h39;
	13'h1DDB: q=8'hBD;
	13'h1DDC: q=8'h0;
	13'h1DDD: q=8'hEB;
	13'h1DDE: q=8'hC6;
	13'h1DDF: q=8'h1;
	13'h1DE0: q=8'hD7;
	13'h1DE1: q=8'h86;
	13'h1DE2: q=8'hBD;
	13'h1DE3: q=8'hEB;
	13'h1DE4: q=8'h1B;
	13'h1DE5: q=8'h7F;
	13'h1DE6: q=8'h0;
	13'h1DE7: q=8'h86;
	13'h1DE8: q=8'hBD;
	13'h1DE9: q=8'hE9;
	13'h1DEA: q=8'hE;
	13'h1DEB: q=8'hEC;
	13'h1DEC: q=8'h2;
	13'h1DED: q=8'hBD;
	13'h1DEE: q=8'hE2;
	13'h1DEF: q=8'h2D;
	13'h1DF0: q=8'hFF;
	13'h1DF1: q=8'h42;
	13'h1DF2: q=8'h71;
	13'h1DF3: q=8'hDE;
	13'h1DF4: q=8'h89;
	13'h1DF5: q=8'hE6;
	13'h1DF6: q=8'h4;
	13'h1DF7: q=8'h58;
	13'h1DF8: q=8'hCB;
	13'h1DF9: q=8'h5;
	13'h1DFA: q=8'h3A;
	13'h1DFB: q=8'hFF;
	13'h1DFC: q=8'h42;
	13'h1DFD: q=8'h6F;
	13'h1DFE: q=8'hBD;
	13'h1DFF: q=8'h0;
	13'h1E00: q=8'hF3;
	13'h1E01: q=8'h27;
	13'h1E02: q=8'hCC;
	13'h1E03: q=8'h7E;
	13'h1E04: q=8'hEA;
	13'h1E05: q=8'h2F;
	13'h1E06: q=8'hBD;
	13'h1E07: q=8'h0;
	13'h1E08: q=8'hEB;
	13'h1E09: q=8'h86;
	13'h1E0A: q=8'h2;
	13'h1E0B: q=8'h8D;
	13'h1E0C: q=8'h82;
	13'h1E0D: q=8'hCE;
	13'h1E0E: q=8'h0;
	13'h1E0F: q=8'h0;
	13'h1E10: q=8'hBD;
	13'h1E11: q=8'h0;
	13'h1E12: q=8'hF3;
	13'h1E13: q=8'h27;
	13'h1E14: q=8'h6;
	13'h1E15: q=8'hBD;
	13'h1E16: q=8'hEA;
	13'h1E17: q=8'h2F;
	13'h1E18: q=8'hBD;
	13'h1E19: q=8'hEF;
	13'h1E1A: q=8'h4C;
	13'h1E1B: q=8'hDF;
	13'h1E1C: q=8'h89;
	13'h1E1D: q=8'hFC;
	13'h1E1E: q=8'h42;
	13'h1E1F: q=8'h6A;
	13'h1E20: q=8'hD3;
	13'h1E21: q=8'h89;
	13'h1E22: q=8'hFD;
	13'h1E23: q=8'h42;
	13'h1E24: q=8'h1F;
	13'h1E25: q=8'hFC;
	13'h1E26: q=8'h42;
	13'h1E27: q=8'h6C;
	13'h1E28: q=8'hD3;
	13'h1E29: q=8'h89;
	13'h1E2A: q=8'h37;
	13'h1E2B: q=8'h36;
	13'h1E2C: q=8'h38;
	13'h1E2D: q=8'h20;
	13'h1E2E: q=8'h99;
	13'h1E2F: q=8'hBD;
	13'h1E30: q=8'hFD;
	13'h1E31: q=8'hA2;
	13'h1E32: q=8'h8D;
	13'h1E33: q=8'h56;
	13'h1E34: q=8'h26;
	13'h1E35: q=8'h9D;
	13'h1E36: q=8'h39;
	13'h1E37: q=8'h96;
	13'h1E38: q=8'hE2;
	13'h1E39: q=8'h4C;
	13'h1E3A: q=8'h26;
	13'h1E3B: q=8'hA;
	13'h1E3C: q=8'hBD;
	13'h1E3D: q=8'hFB;
	13'h1E3E: q=8'hD4;
	13'h1E3F: q=8'h86;
	13'h1E40: q=8'h53;
	13'h1E41: q=8'h8D;
	13'h1E42: q=8'h3E;
	13'h1E43: q=8'hBD;
	13'h1E44: q=8'hE7;
	13'h1E45: q=8'hB9;
	13'h1E46: q=8'h8D;
	13'h1E47: q=8'h62;
	13'h1E48: q=8'hBA;
	13'h1E49: q=8'h42;
	13'h1E4A: q=8'h75;
	13'h1E4B: q=8'h26;
	13'h1E4C: q=8'h33;
	13'h1E4D: q=8'h5F;
	13'h1E4E: q=8'h37;
	13'h1E4F: q=8'hCE;
	13'h1E50: q=8'h42;
	13'h1E51: q=8'h5F;
	13'h1E52: q=8'h3A;
	13'h1E53: q=8'hA6;
	13'h1E54: q=8'h0;
	13'h1E55: q=8'hDE;
	13'h1E56: q=8'hE2;
	13'h1E57: q=8'h8;
	13'h1E58: q=8'h26;
	13'h1E59: q=8'h2;
	13'h1E5A: q=8'h8D;
	13'h1E5B: q=8'h25;
	13'h1E5C: q=8'hCE;
	13'h1E5D: q=8'h42;
	13'h1E5E: q=8'h57;
	13'h1E5F: q=8'h3A;
	13'h1E60: q=8'hA0;
	13'h1E61: q=8'h0;
	13'h1E62: q=8'h30;
	13'h1E63: q=8'hAA;
	13'h1E64: q=8'h0;
	13'h1E65: q=8'hA7;
	13'h1E66: q=8'h0;
	13'h1E67: q=8'h5C;
	13'h1E68: q=8'hC1;
	13'h1E69: q=8'h8;
	13'h1E6A: q=8'h26;
	13'h1E6B: q=8'hE3;
	13'h1E6C: q=8'h32;
	13'h1E6D: q=8'h4D;
	13'h1E6E: q=8'h27;
	13'h1E6F: q=8'hB;
	13'h1E70: q=8'h7D;
	13'h1E71: q=8'h42;
	13'h1E72: q=8'h56;
	13'h1E73: q=8'h27;
	13'h1E74: q=8'h6;
	13'h1E75: q=8'h8D;
	13'h1E76: q=8'h10;
	13'h1E77: q=8'h26;
	13'h1E78: q=8'h7;
	13'h1E79: q=8'h20;
	13'h1E7A: q=8'hBC;
	13'h1E7B: q=8'h86;
	13'h1E7C: q=8'h46;
	13'h1E7D: q=8'h8D;
	13'h1E7E: q=8'h22;
	13'h1E7F: q=8'h4F;
	13'h1E80: q=8'h39;
	13'h1E81: q=8'h7F;
	13'h1E82: q=8'h0;
	13'h1E83: q=8'hE8;
	13'h1E84: q=8'h7E;
	13'h1E85: q=8'hF9;
	13'h1E86: q=8'hC6;
	13'h1E87: q=8'hBD;
	13'h1E88: q=8'hFF;
	13'h1E89: q=8'h4E;
	13'h1E8A: q=8'h86;
	13'h1E8B: q=8'hFF;
	13'h1E8C: q=8'h16;
	13'h1E8D: q=8'h8D;
	13'h1E8E: q=8'h2A;
	13'h1E8F: q=8'h26;
	13'h1E90: q=8'h7;
	13'h1E91: q=8'hB6;
	13'h1E92: q=8'h42;
	13'h1E93: q=8'h75;
	13'h1E94: q=8'h40;
	13'h1E95: q=8'h2B;
	13'h1E96: q=8'hF3;
	13'h1E97: q=8'h4A;
	13'h1E98: q=8'hB7;
	13'h1E99: q=8'h42;
	13'h1E9A: q=8'h7B;
	13'h1E9B: q=8'h39;
	13'h1E9C: q=8'hB6;
	13'h1E9D: q=8'h40;
	13'h1E9E: q=8'h0;
	13'h1E9F: q=8'h88;
	13'h1EA0: q=8'h40;
	13'h1EA1: q=8'hD6;
	13'h1EA2: q=8'hE2;
	13'h1EA3: q=8'h5C;
	13'h1EA4: q=8'h26;
	13'h1EA5: q=8'h3;
	13'h1EA6: q=8'hB7;
	13'h1EA7: q=8'h40;
	13'h1EA8: q=8'h0;
	13'h1EA9: q=8'h39;
	13'h1EAA: q=8'hBD;
	13'h1EAB: q=8'hFF;
	13'h1EAC: q=8'h4E;
	13'h1EAD: q=8'hCE;
	13'h1EAE: q=8'h42;
	13'h1EAF: q=8'h5F;
	13'h1EB0: q=8'hFF;
	13'h1EB1: q=8'h42;
	13'h1EB2: q=8'h78;
	13'h1EB3: q=8'h86;
	13'h1EB4: q=8'hF;
	13'h1EB5: q=8'h8C;
	13'h1EB6: q=8'h86;
	13'h1EB7: q=8'hFF;
	13'h1EB8: q=8'h5F;
	13'h1EB9: q=8'h36;
	13'h1EBA: q=8'hF7;
	13'h1EBB: q=8'h42;
	13'h1EBC: q=8'h73;
	13'h1EBD: q=8'h1;
	13'h1EBE: q=8'hF;
	13'h1EBF: q=8'h8D;
	13'h1EC0: q=8'hDB;
	13'h1EC1: q=8'hFE;
	13'h1EC2: q=8'h42;
	13'h1EC3: q=8'h78;
	13'h1EC4: q=8'h4F;
	13'h1EC5: q=8'h8D;
	13'h1EC6: q=8'h5B;
	13'h1EC7: q=8'h46;
	13'h1EC8: q=8'h81;
	13'h1EC9: q=8'h3C;
	13'h1ECA: q=8'h26;
	13'h1ECB: q=8'hF9;
	13'h1ECC: q=8'h8D;
	13'h1ECD: q=8'h46;
	13'h1ECE: q=8'hB7;
	13'h1ECF: q=8'h42;
	13'h1ED0: q=8'h75;
	13'h1ED1: q=8'h8D;
	13'h1ED2: q=8'h41;
	13'h1ED3: q=8'hB7;
	13'h1ED4: q=8'h42;
	13'h1ED5: q=8'h76;
	13'h1ED6: q=8'h33;
	13'h1ED7: q=8'h11;
	13'h1ED8: q=8'h22;
	13'h1ED9: q=8'h31;
	13'h1EDA: q=8'hBB;
	13'h1EDB: q=8'h42;
	13'h1EDC: q=8'h75;
	13'h1EDD: q=8'hB7;
	13'h1EDE: q=8'h42;
	13'h1EDF: q=8'h7A;
	13'h1EE0: q=8'hB6;
	13'h1EE1: q=8'h42;
	13'h1EE2: q=8'h76;
	13'h1EE3: q=8'hB7;
	13'h1EE4: q=8'h42;
	13'h1EE5: q=8'h7B;
	13'h1EE6: q=8'h27;
	13'h1EE7: q=8'h19;
	13'h1EE8: q=8'h8D;
	13'h1EE9: q=8'h2A;
	13'h1EEA: q=8'h7D;
	13'h1EEB: q=8'h42;
	13'h1EEC: q=8'h73;
	13'h1EED: q=8'h26;
	13'h1EEE: q=8'h7;
	13'h1EEF: q=8'hA7;
	13'h1EF0: q=8'h0;
	13'h1EF1: q=8'hA1;
	13'h1EF2: q=8'h0;
	13'h1EF3: q=8'h26;
	13'h1EF4: q=8'h19;
	13'h1EF5: q=8'h8;
	13'h1EF6: q=8'hBB;
	13'h1EF7: q=8'h42;
	13'h1EF8: q=8'h7A;
	13'h1EF9: q=8'hB7;
	13'h1EFA: q=8'h42;
	13'h1EFB: q=8'h7A;
	13'h1EFC: q=8'h7A;
	13'h1EFD: q=8'h42;
	13'h1EFE: q=8'h7B;
	13'h1EFF: q=8'h26;
	13'h1F00: q=8'hE7;
	13'h1F01: q=8'h8D;
	13'h1F02: q=8'h11;
	13'h1F03: q=8'hB0;
	13'h1F04: q=8'h42;
	13'h1F05: q=8'h7A;
	13'h1F06: q=8'h27;
	13'h1F07: q=8'h8;
	13'h1F08: q=8'h86;
	13'h1F09: q=8'h1;
	13'h1F0A: q=8'h8C;
	13'h1F0B: q=8'h86;
	13'h1F0C: q=8'h3;
	13'h1F0D: q=8'h8C;
	13'h1F0E: q=8'h86;
	13'h1F0F: q=8'h2;
	13'h1F10: q=8'hB7;
	13'h1F11: q=8'h42;
	13'h1F12: q=8'h7B;
	13'h1F13: q=8'h39;
	13'h1F14: q=8'h86;
	13'h1F15: q=8'h8;
	13'h1F16: q=8'hB7;
	13'h1F17: q=8'h42;
	13'h1F18: q=8'h7C;
	13'h1F19: q=8'h8D;
	13'h1F1A: q=8'h7;
	13'h1F1B: q=8'h46;
	13'h1F1C: q=8'h7A;
	13'h1F1D: q=8'h42;
	13'h1F1E: q=8'h7C;
	13'h1F1F: q=8'h26;
	13'h1F20: q=8'hF8;
	13'h1F21: q=8'h39;
	13'h1F22: q=8'h8D;
	13'h1F23: q=8'h8;
	13'h1F24: q=8'hF6;
	13'h1F25: q=8'h42;
	13'h1F26: q=8'h7D;
	13'h1F27: q=8'h5A;
	13'h1F28: q=8'hF1;
	13'h1F29: q=8'h42;
	13'h1F2A: q=8'h2C;
	13'h1F2B: q=8'h39;
	13'h1F2C: q=8'h7F;
	13'h1F2D: q=8'h42;
	13'h1F2E: q=8'h7D;
	13'h1F2F: q=8'h7D;
	13'h1F30: q=8'h42;
	13'h1F31: q=8'h7E;
	13'h1F32: q=8'h26;
	13'h1F33: q=8'h11;
	13'h1F34: q=8'h8D;
	13'h1F35: q=8'h7;
	13'h1F36: q=8'h26;
	13'h1F37: q=8'hFC;
	13'h1F38: q=8'h8D;
	13'h1F39: q=8'h3;
	13'h1F3A: q=8'h27;
	13'h1F3B: q=8'hFC;
	13'h1F3C: q=8'h39;
	13'h1F3D: q=8'h7C;
	13'h1F3E: q=8'h42;
	13'h1F3F: q=8'h7D;
	13'h1F40: q=8'hD6;
	13'h1F41: q=8'h3;
	13'h1F42: q=8'hC4;
	13'h1F43: q=8'h10;
	13'h1F44: q=8'h39;
	13'h1F45: q=8'h8D;
	13'h1F46: q=8'hF6;
	13'h1F47: q=8'h27;
	13'h1F48: q=8'hFC;
	13'h1F49: q=8'h8D;
	13'h1F4A: q=8'hF2;
	13'h1F4B: q=8'h26;
	13'h1F4C: q=8'hFC;
	13'h1F4D: q=8'h39;
	13'h1F4E: q=8'h1;
	13'h1F4F: q=8'hF;
	13'h1F50: q=8'h7F;
	13'h1F51: q=8'h42;
	13'h1F52: q=8'h7C;
	13'h1F53: q=8'h8D;
	13'h1F54: q=8'hDF;
	13'h1F55: q=8'h8D;
	13'h1F56: q=8'h2D;
	13'h1F57: q=8'h22;
	13'h1F58: q=8'h12;
	13'h1F59: q=8'h8D;
	13'h1F5A: q=8'h22;
	13'h1F5B: q=8'h25;
	13'h1F5C: q=8'h12;
	13'h1F5D: q=8'h7A;
	13'h1F5E: q=8'h42;
	13'h1F5F: q=8'h7C;
	13'h1F60: q=8'hB6;
	13'h1F61: q=8'h42;
	13'h1F62: q=8'h7C;
	13'h1F63: q=8'h81;
	13'h1F64: q=8'hA0;
	13'h1F65: q=8'h26;
	13'h1F66: q=8'hEC;
	13'h1F67: q=8'hB7;
	13'h1F68: q=8'h42;
	13'h1F69: q=8'h7E;
	13'h1F6A: q=8'h39;
	13'h1F6B: q=8'h8D;
	13'h1F6C: q=8'h10;
	13'h1F6D: q=8'h22;
	13'h1F6E: q=8'hE6;
	13'h1F6F: q=8'h8D;
	13'h1F70: q=8'h13;
	13'h1F71: q=8'h25;
	13'h1F72: q=8'hE6;
	13'h1F73: q=8'h7C;
	13'h1F74: q=8'h42;
	13'h1F75: q=8'h7C;
	13'h1F76: q=8'hB6;
	13'h1F77: q=8'h42;
	13'h1F78: q=8'h7C;
	13'h1F79: q=8'h80;
	13'h1F7A: q=8'h60;
	13'h1F7B: q=8'h20;
	13'h1F7C: q=8'hE8;
	13'h1F7D: q=8'h7F;
	13'h1F7E: q=8'h42;
	13'h1F7F: q=8'h7D;
	13'h1F80: q=8'h8D;
	13'h1F81: q=8'hB6;
	13'h1F82: q=8'h20;
	13'h1F83: q=8'h5;
	13'h1F84: q=8'h7F;
	13'h1F85: q=8'h42;
	13'h1F86: q=8'h7D;
	13'h1F87: q=8'h8D;
	13'h1F88: q=8'hC0;
	13'h1F89: q=8'hF6;
	13'h1F8A: q=8'h42;
	13'h1F8B: q=8'h7D;
	13'h1F8C: q=8'hF1;
	13'h1F8D: q=8'h42;
	13'h1F8E: q=8'h2D;
	13'h1F8F: q=8'h22;
	13'h1F90: q=8'h4;
	13'h1F91: q=8'hF1;
	13'h1F92: q=8'h42;
	13'h1F93: q=8'h2E;
	13'h1F94: q=8'h39;
	13'h1F95: q=8'h7F;
	13'h1F96: q=8'h42;
	13'h1F97: q=8'h7C;
	13'h1F98: q=8'h39;
	13'h1F99: q=8'hBD;
	13'h1F9A: q=8'hEA;
	13'h1F9B: q=8'h2F;
	13'h1F9C: q=8'hBD;
	13'h1F9D: q=8'hEF;
	13'h1F9E: q=8'hD;
	13'h1F9F: q=8'h5D;
	13'h1FA0: q=8'h26;
	13'h1FA1: q=8'h2F;
	13'h1FA2: q=8'h7E;
	13'h1FA3: q=8'hEC;
	13'h1FA4: q=8'h2E;
	13'h1FA5: q=8'h8D;
	13'h1FA6: q=8'hF5;
	13'h1FA7: q=8'h37;
	13'h1FA8: q=8'h8D;
	13'h1FA9: q=8'hEF;
	13'h1FAA: q=8'h32;
	13'h1FAB: q=8'h36;
	13'h1FAC: q=8'h37;
	13'h1FAD: q=8'h4F;
	13'h1FAE: q=8'hDE;
	13'h1FAF: q=8'h9;
	13'h1FB0: q=8'hD6;
	13'h1FB1: q=8'h8;
	13'h1FB2: q=8'hDF;
	13'h1FB3: q=8'hB;
	13'h1FB4: q=8'h88;
	13'h1FB5: q=8'h80;
	13'h1FB6: q=8'hB7;
	13'h1FB7: q=8'hBF;
	13'h1FB8: q=8'hFF;
	13'h1FB9: q=8'h30;
	13'h1FBA: q=8'hE6;
	13'h1FBB: q=8'h1;
	13'h1FBC: q=8'h8;
	13'h1FBD: q=8'h8;
	13'h1FBE: q=8'h5C;
	13'h1FBF: q=8'h26;
	13'h1FC0: q=8'hFB;
	13'h1FC1: q=8'hD6;
	13'h1FC2: q=8'h8;
	13'h1FC3: q=8'hC4;
	13'h1FC4: q=8'h40;
	13'h1FC5: q=8'h27;
	13'h1FC6: q=8'hED;
	13'h1FC7: q=8'h30;
	13'h1FC8: q=8'h6A;
	13'h1FC9: q=8'h0;
	13'h1FCA: q=8'h26;
	13'h1FCB: q=8'hE2;
	13'h1FCC: q=8'h4F;
	13'h1FCD: q=8'hB7;
	13'h1FCE: q=8'hBF;
	13'h1FCF: q=8'hFF;
	13'h1FD0: q=8'h38;
	13'h1FD1: q=8'h39;
	13'h1FD2: q=8'h6E;
	13'h1FD3: q=8'h69;
	13'h1FD4: q=8'h6C;
	13'h1FD5: q=8'h72;
	13'h1FD6: q=8'h65;
	13'h1FD7: q=8'h62;
	13'h1FD8: q=8'h6D;
	13'h1FD9: q=8'h61;
	13'h1FDA: q=8'h68;
	13'h1FDB: q=8'h43;
	13'h1FDC: q=8'hF8;
	13'h1FDD: q=8'h83;
	13'h1FDE: q=8'hF9;
	13'h1FDF: q=8'hC6;
	13'h1FE0: q=8'hFF;
	13'h1FE1: q=8'h4E;
	13'h1FE2: q=8'hFE;
	13'h1FE3: q=8'hB9;
	13'h1FE4: q=8'hFC;
	13'h1FE5: q=8'hC0;
	13'h1FE6: q=8'hFF;
	13'h1FE7: q=8'hAB;
	13'h1FE8: q=8'hFC;
	13'h1FE9: q=8'hB7;
	13'h1FEA: q=8'hEC;
	13'h1FEB: q=8'hE3;
	13'h1FEC: q=8'hEB;
	13'h1FED: q=8'hC7;
	13'h1FEE: q=8'h0;
	13'h1FEF: q=8'hC9;
	13'h1FF0: q=8'h42;
	13'h1FF1: q=8'h0;
	13'h1FF2: q=8'h42;
	13'h1FF3: q=8'h3;
	13'h1FF4: q=8'h42;
	13'h1FF5: q=8'h6;
	13'h1FF6: q=8'h42;
	13'h1FF7: q=8'h9;
	13'h1FF8: q=8'h42;
	13'h1FF9: q=8'hC;
	13'h1FFA: q=8'h42;
	13'h1FFB: q=8'hF;
	13'h1FFC: q=8'h42;
	13'h1FFD: q=8'h12;
	13'h1FFE: q=8'hF7;
	13'h1FFF: q=8'h2E;
endcase
end
assign dout = ~cs ? q : 8'd0;
endmodule
